From stdpp Require Import prelude.
From Coq Require Import Streams.
From VLSM.Lib Require Import Preamble ListExtras StreamExtras.

(** * VLSM Basics

This module provides basic VLSM infrastructure.
*)

(** ** VLSM definition

*** The type of a VLSM

The type of a VLSM is a triple consisting of the underlying types of
messages, states, and labels.

In Coq it is defined as a Class taking <<message>> as parameter and having
[state] and [label] as fields.  <<message>> is a parameter to allow it to be
easily shared by multiple VLSMs during composition.
*)

Class VLSMType (message : Type) :=
  { state : Type
  ; label : Type
  }.

(** *** The signature of a VLSM

Although the VLSM definition does not single out the notion of a VLSM
signature, we find it convenient to extract it as the [VLSMSign] class.

The [VLSMSign] class is parameterized by a [VLSMType] and defines properties
for initial states ([initial_state_prop]) and initial messages
([initial_message_prop]), from which we can immediately define the dependent
types [initial_state] (as [state]s having the [initial_state_prop]erty) and
[intial_message] (as <<message>>s having the [initial_message_prop]erty).

Additionally, [VLSMSign] requires the identification of an [initial_state] [s0],
a <<message>> [m0], and a [label] [l0] to ensure the non-emptiness of the
corresponding sets.
*)

  Class VLSMSign {message : Type} (vtype : VLSMType message) :=
    { initial_state_prop : state -> Prop
    ; initial_state := { s : state | initial_state_prop s }
    ; initial_message_prop : message -> Prop
    ; initial_message := { m : message | initial_message_prop m }
    ; s0 : Inhabited initial_state
    }.

  Definition option_initial_message_prop
    {message : Type} {vtype : VLSMType message} {sign : VLSMSign vtype}
    : option message -> Prop := from_option initial_message_prop True.

  Definition VLSMSign_pre_loaded_with_messages
    {message : Type} {vtype : VLSMType message} (sign : VLSMSign vtype)
    (initial : message -> Prop)
    : VLSMSign vtype
    :=
    {| initial_state_prop := @initial_state_prop _ _ sign
    ; initial_message_prop := fun m => @initial_message_prop _ _ sign  m \/ initial m
    ; s0 := @s0 _ _ sign
    |}.

  Definition decidable_initial_messages_prop
    {message : Type} {vtype : VLSMType message} (sign : VLSMSign vtype)
    := forall m, Decision (initial_message_prop m).

(** *** VLSM class definition

Given a [VLSMSign]nature, a [VLSM] is defined by providing a [transition]
function and a [valid]ity condition.
*)

  Class VLSMClass {message : Type} {vtype : VLSMType message} (lsm : VLSMSign vtype) :=
    { transition : label -> state * option message -> state * option message
    ; valid : label -> state * option message -> Prop
    }.

  Definition VLSMClass_pre_loaded_with_messages
    {message : Type} {vtype : VLSMType message} {lsm : VLSMSign vtype} (vlsm : VLSMClass lsm)
    (initial : message -> Prop)
    : VLSMClass (VLSMSign_pre_loaded_with_messages lsm initial)
    :=
    {| transition := @transition _ _ _ vlsm
     ; valid := @valid _ _ _ vlsm
    |}.

  (** For technical reasons, e.g., the need to easily talk about VLSMs over
  the same set of messages and about VLSMs of the same type (over the same
  set of messages, labels and states), the VLSM definition is split into
  three parts, [VLSM_Type], [VLSM_Sign], and [VLSMClass], which are
  packaged together by the following definition.
  *)
  Definition VLSM (message : Type) :=
    sigT (fun T : VLSMType message =>
      sigT (fun S : VLSMSign T => VLSMClass S)).

  Definition mk_vlsm
    {message : Type}
    {T : VLSMType message}
    {S : VLSMSign T}
    (M : VLSMClass S)
    : VLSM message
    := existT T (existT S M).

  Definition pre_loaded_vlsm
    {message : Type}
    (X : VLSM message)
    (initial : message -> Prop)
    : VLSM message
    :=
    let M := projT2 (projT2 X) in
    let M' := VLSMClass_pre_loaded_with_messages M initial in
    mk_vlsm M'.

Section Traces.

  Context
    {message : Type}
    {T : VLSMType message}
    .

(** ** Traces

We introduce the concept of a trace to formalize an execution of the protocol.
It is abstracted as a pair <<(start, steps)>> where <<start>> is a state
and <<steps>> is a tuple of objects which fully describe the transitions
underwent during execution. Notably, <<steps>> might be infinite.

In Coq, we can define these objects (which we name [transition_item]s) as consisting of:
- the [label] [l]
- the (optional) [input] <<message>>
- the [destination] [state] of the transition
- the (optional) [output] <<message>> generated by the transition
*)

  Record transition_item :=
    {   l : label
        ;   input : option message
        ;   destination : state
        ;   output : option message
    }.

    Definition field_selector
               (field: transition_item -> option message) :
      (message -> transition_item -> Prop) :=
      fun m item => field item = Some m.

    Definition item_sends_or_receives:
      message -> transition_item -> Prop :=
      fun m item => input item = Some m \/ output item = Some m.

    Definition trace_has_message
      (message_selector : message -> transition_item -> Prop)
      (msg : message)
      (tr : list transition_item)
      : Prop
      := List.Exists (message_selector msg) tr.

    Lemma trace_has_message_prefix
      (message_selector : message -> transition_item -> Prop)
      (msg : message)
      (prefix suffix : list transition_item)
      : trace_has_message message_selector msg prefix ->
        trace_has_message message_selector msg (prefix ++ suffix).
    Proof.
      intro Hprefix.
      apply Exists_app. left. assumption.
    Qed.

    Lemma trace_has_message_observed_iff m tr
      (Hobserved : trace_has_message item_sends_or_receives m tr)
      : trace_has_message (field_selector input) m tr \/ trace_has_message (field_selector output) m tr.
    Proof.
      unfold trace_has_message in *. rewrite !Exists_exists in *.
      destruct Hobserved as [item [Hitem [Hm|Hm]]]
      ; [left|right]; exists item; split; assumption.
    Qed.

    (** Defines a message received but not sent by within the trace. *)
    Definition trace_received_not_sent_before_or_after
      (tr : list transition_item)
      (m : message)
      : Prop
      := trace_has_message (field_selector input) m tr /\
         ~trace_has_message (field_selector output) m tr.

    (** States that a property holds for all messages received but not sent by a trace. *)
    Definition trace_received_not_sent_before_or_after_invariant
      (tr : list transition_item)
      (P : message -> Prop)
      : Prop
      := forall m, trace_received_not_sent_before_or_after tr m -> P m.

  (** [proto_run] is used for an alternative definition of [valid_state_message_prop], which
  takes into account transitions. See 'vlsm_run_prop'.
  *)
  Record proto_run : Type := mk_proto_run
    { start : state
      ; transitions : list transition_item
      ; final : state * option message
    }.

  Inductive Trace : Type :=
  | Finite : state -> list transition_item -> Trace
  | Infinite : state -> Stream transition_item -> Trace.

  Definition trace_first (tr : Trace) : state :=
    match tr with
    | Finite s _ => s
    | Infinite s _ => s
    end.

  Definition finite_trace_last
    (si : state) (tr : list transition_item) : state :=
    List.last (List.map destination tr) si.

  Definition finite_trace_last_output
    (tr : list transition_item) : option message :=
    List.last (List.map output tr) None.

  Definition finite_trace_nth
    (si : state) (tr : list transition_item)
    : nat -> option state :=
  nth_error (si :: List.map destination tr).

  Definition trace_last (tr : Trace) : option state
    :=
      match tr with
      | Finite s ls => Some (finite_trace_last s ls)
      | Infinite _ _ => None
      end.

(**
Next function extract the nth state of a trace, where the sequence of
states of a trace is obtained by appending the all destination
states in the transition list/stream to the initial state of the trace.
*)
  Definition trace_nth (tr : Trace)
    : nat -> option state :=
    fun (n : nat) =>
      match tr with
      | Finite s ls => finite_trace_nth s ls n
      | Infinite s st => Some (Str_nth n (Cons s (Streams.map destination st)))
      end.

End Traces.

Arguments transition_item {message} {T} , {message} T.
Arguments field_selector {_} {T} _ msg item / .
Arguments item_sends_or_receives {_} {_} msg item /.

Section TraceLemmas.

  Context
    [message : Type]
    [T : VLSMType message]
    .

  Lemma last_error_destination_last
    (tr : list transition_item)
    (s : state)
    (Hlast : option_map destination (last_error tr) = Some s)
    (default : state)
    : finite_trace_last default tr  = s.
  Proof.
    unfold option_map in Hlast.
    destruct (last_error tr) eqn : eq; try discriminate Hlast.
    inversion Hlast.
    unfold last_error in eq.
    destruct tr; try discriminate eq.
    inversion eq.
    unfold finite_trace_last.
    rewrite last_map. reflexivity.
  Qed.

  Lemma finite_trace_last_cons
    s x tl:
    finite_trace_last s (x::tl) = finite_trace_last (destination x) tl.
  Proof.
    unfold finite_trace_last. rewrite map_cons, unroll_last. reflexivity.
  Qed.

  Lemma finite_trace_last_nil
    s:
    finite_trace_last s [] = s.
  Proof. reflexivity. Qed.

  Lemma finite_trace_last_app
    s t1 t2:
    finite_trace_last s (t1 ++ t2) = finite_trace_last (finite_trace_last s t1) t2.
  Proof.
    unfold finite_trace_last.
    rewrite map_app, last_app.
    reflexivity.
  Qed.

  Lemma finite_trace_last_is_last
    s x tl:
    finite_trace_last s (tl++[x]) = destination x.
  Proof.
    unfold finite_trace_last.
    rewrite map_app.
    simpl.
    rewrite last_is_last.
    reflexivity.
  Qed.

  Lemma finite_trace_last_output_is_last
    x tl:
    finite_trace_last_output (tl++[x]) = output x.
  Proof.
    unfold finite_trace_last_output.
    rewrite map_app.
    simpl.
    rewrite last_is_last.
    reflexivity.
  Qed.

  Lemma finite_trace_nth_first
    (si : state) (tr : list transition_item):
    finite_trace_nth si tr 0 = Some si.
  Proof.
    reflexivity.
  Qed.

  Lemma finite_trace_nth_last
    (si : state) (tr : list transition_item):
    finite_trace_nth si tr (length tr) = Some (finite_trace_last si tr).
  Proof.
    unfold finite_trace_nth, finite_trace_last.
    destruct tr;[reflexivity|].
    cbn [nth_error length].
    apply nth_error_last.
    rewrite map_length.
    reflexivity.
  Qed.

  Lemma finite_trace_nth_app1
    (si : state) (t1 t2 : list transition_item) n:
    n <= length t1 ->
    finite_trace_nth si (t1++t2) n = finite_trace_nth si t1 n.
  Proof.
    intro H.
    unfold finite_trace_nth.
    rewrite map_app, app_comm_cons.
    apply nth_error_app1.
    simpl. rewrite map_length.
    auto with arith.
  Qed.

  Lemma finite_trace_nth_app2
    (si : state) (t1 t2 : list transition_item) n:
    length t1 <= n ->
    finite_trace_nth si (t1++t2) n = finite_trace_nth (finite_trace_last si t1) t2 (n - length t1).
  Proof.
    intro H.
    apply Compare_dec.le_lt_eq_dec in H.
    destruct H as [H |<-].
    - unfold finite_trace_nth.
      rewrite map_app, app_comm_cons.
      rewrite nth_error_app2;simpl length;rewrite map_length;[|solve[auto with arith]].
      destruct n;[exfalso;lia|].
      replace (S n -length t1) with (S (n - length t1)) by lia.
      reflexivity.
    - rewrite finite_trace_nth_app1, finite_trace_nth_last by reflexivity.
      rewrite PeanoNat.Nat.sub_diag, finite_trace_nth_first.
      reflexivity.
  Qed.

  Lemma finite_trace_nth_length
    (si : state) (tr : list transition_item) n s:
    finite_trace_nth si tr n = Some s ->
    n <= length tr.
  Proof.
    intros H.
    apply nth_error_length in H.
    simpl in H.
    rewrite map_length in H.
    apply le_S_n in H.
    assumption.
  Qed.

  Lemma finite_trace_last_prefix
    (s: state) (tr: list transition_item) n nth:
    finite_trace_nth s tr n = Some nth ->
    finite_trace_last s (list_prefix tr n) = nth.
  Proof.
    unfold finite_trace_nth, finite_trace_last.
    rewrite list_prefix_map.
    generalize (List.map destination tr); intro l; clear tr.
    destruct n.
    - simpl. intros [=<-]. destruct l;reflexivity.
    - simpl. intro H. symmetry. revert H s.
      apply list_prefix_nth_last.
  Qed.

  Lemma finite_trace_last_suffix
    (s: state) (tr: list transition_item) n:
    n < length tr ->
    finite_trace_last s (list_suffix tr n) = finite_trace_last s tr.
  Proof.
    intros H.
    unfold finite_trace_last.
    rewrite list_suffix_map.
    apply list_suffix_last.
    rewrite map_length.
    assumption.
  Qed.

  Lemma unlock_finite_trace_last s tr:
    finite_trace_last s tr = List.last (List.map destination tr) s.
  Proof.
    reflexivity.
  Qed.
  Opaque finite_trace_last.

End TraceLemmas.

Section vlsm_projections.

  Context
    {message : Type}
    (vlsm : VLSM message)
    .

(**
Given a [VLSM], it is convenient to be able to retrieve its V[VLSMSign]nature
or [VLSMType]. Functions [sign] and [type] below achieve this precise purpose.
*)

  Definition type := projT1 vlsm.
  Definition sign := projT1 (projT2 vlsm).
  Definition machine := projT2 (projT2 vlsm).
  Definition vstate := @state _ type.
  Definition vlabel := @label _ type.
  Definition vinitial_state_prop := @initial_state_prop _ _ sign.
  Definition vinitial_state := @initial_state _ _ sign.
  Definition vinitial_message_prop := @initial_message_prop _ _ sign.
  Definition voption_initial_message_prop := @option_initial_message_prop _ _ sign.
  Definition vinitial_message := @initial_message _ _ sign.
  Definition vs0 := @inhabitant _ (@s0 _ _ sign).
  Definition vdecidable_initial_messages_prop := @decidable_initial_messages_prop _ _ sign.
  Definition vtransition := @transition _ _ _ machine.
  Definition vvalid := @valid _ _ _ machine.
  Definition vtransition_item := @transition_item _ type.
  Definition vTrace := @Trace _ type.
  Definition vproto_run := @proto_run _ type.

End vlsm_projections.

Ltac unfold_vtransition H := (unfold vtransition in H; simpl in H).

Lemma mk_vlsm_machine
  {message : Type}
  (X : VLSM message)
  : mk_vlsm (machine X) = X.
Proof.
  destruct X as (T, (S, M)). reflexivity.
Qed.

  Section VLSM.

(**
In this section we assume a fixed [VLSM].
*)

    Context
      {message : Type}
      (X : VLSM message)
      (TypeX := type X)
      (SignX := sign X)
      (MachineX := machine X)
      .

Existing Instance TypeX.
Existing Instance SignX.
Existing Instance MachineX.

(** *** Valid states and messages

We further characterize certain objects as being _valid_, which means they can
be witnessed or experienced during executions of the protocol. For example,
a message is a [valid_message] if there exists an execution of the protocol
in which it is produced.

We choose here to define valid states and messages together as the
[valid_state_message_prop]erty, inductively defined over the
[state * option message] product type,
as this definition avoids the need of using a mutually recursive definition.

The inductive definition has three cases:
- if <<s>> is a [state] with the [initial_state_prop]erty, then <<(s, None)>>
  has the [valid_state_message_prop]erty;
- if <<m>> is a <<message>> with the [initial_message_prop]erty,
  then <<(>>[s0, Some]<< m)>> has the [valid_state_message_prop]erty;
- for all [state]s <<s>>, [option]al <<message>> <<om>>, and [label] <<l>>:

  - if there is an (optional) <<message>> <<_om>> such that <<(s, _om)>>
    has the [valid_state_message_prop]erty;

  - and if there is a [state] <<_s>> such that <<(_s, om)>> has the
    [valid_state_message_prop]erty;

  - and if <<l>> [valid] <<(s, om)>>,

  - then [transition] <<l (s, om)>> has the [valid_state_message_prop]erty.
*)

    Inductive valid_state_message_prop : state -> option message -> Prop :=
    | valid_initial_state_message
        (s : state)
        (Hs : initial_state_prop s)
        (om : option message)
        (Hom : option_initial_message_prop om)
      : valid_state_message_prop s om
    | valid_generated_state_message
        (s : state)
        (_om : option message)
        (Hps : valid_state_message_prop s _om)
        (_s : state)
        (om : option message)
        (Hpm : valid_state_message_prop _s om)
        (l : label)
        (Hv : valid l (s, om))
        s' om'
        (Ht : transition l (s, om) = (s', om'))
      : valid_state_message_prop s' om'.

    Definition valid_initial_state
      [s:state] (Hs: initial_state_prop s)
      : valid_state_message_prop s None
      := valid_initial_state_message s Hs None I.

(**

The [valid_state_prop]erty and the [valid_message_prop]erty are now
definable as simple projections of the above definition.

Moreover, we use these derived properties to define the corresponding
dependent types [valid_state] and [valid_message].

*)

    Definition valid_state_prop (s : state) :=
      exists om : option message, valid_state_message_prop s om.

    Definition valid_message_prop (m : message) :=
      exists s : state, valid_state_message_prop s (Some m).

    Definition valid_state : Type :=
      { s : state | valid_state_prop s }.

    Definition valid_message : Type :=
      { m : message | valid_message_prop m }.

    Lemma initial_state_is_valid
      (s : state)
      (Hinitial : initial_state_prop s) :
      valid_state_prop s.
    Proof.
      exists None.
      apply valid_initial_state_message.
      assumption.
      exact I.
    Qed.

    Lemma initial_message_is_valid
      (m : message)
      (Hinitial : initial_message_prop m) :
      valid_message_prop m.
    Proof.
      exists (proj1_sig (vs0 X)).
      apply valid_initial_state_message.
      apply proj2_sig.
      assumption.
    Qed.

(**
As often times we work with optional valid messages, it is convenient
to define a valid message property for optional messages:
*)

    Definition option_valid_message_prop (om : option message) :=
      exists s : state, valid_state_message_prop s om.

    Lemma option_valid_message_None
      : option_valid_message_prop None.
    Proof.
      exists (proj1_sig (vs0 X)).
      apply valid_initial_state_message.
      apply proj2_sig.
      exact I.
    Qed.

    Lemma option_valid_message_Some
      (m : message)
      (Hpm : valid_message_prop m)
      : option_valid_message_prop (Some m).
    Proof.
      destruct Hpm as [s Hpm]. exists s. assumption.
    Qed.

    Lemma option_initial_message_is_valid
      (om : option message)
      (Hinitial : option_initial_message_prop om) :
      option_valid_message_prop om.
    Proof.
      destruct om;
      [apply option_valid_message_Some
      |apply option_valid_message_None].
      apply initial_message_is_valid;assumption.
    Qed.

(** *** Input validity and input valid transitions

To specify that a particular (input of a) transition can actually be
encountered as part of a protocol execution, we define the notions of
[input_valid]ity and [input_valid_transition].

Input validity requires that the [valid] predicate holds for the
given inputs and that they have a [valid_state] and a [valid_message].
*)
    Definition input_valid
               (l : label)
               (som : state * option message)
      : Prop
      :=
      let (s, om) := som in
         valid_state_prop s
      /\ option_valid_message_prop om
      /\ valid l (s,om).

(** Input valid transitions are transitions with [input_valid] inputs. *)
    Definition input_valid_transition
      (l : label)
      (som : state * option message)
      (som' : state * option message)
      :=
      input_valid l som
      /\  transition l som = som'.

    Definition input_valid_transition_item
      (s : state)
      (item : transition_item)
      :=
      input_valid_transition (l item) (s, input item) (destination item, output item).

    Definition input_valid_transition_preserving
      (R : state -> state -> Prop)
      : Prop
      :=
      forall
        (s1 s2 : state)
        (l : label)
        (om1 om2 : option message)
        (Hvalid_transition: input_valid_transition l (s1, om1) (s2, om2)),
        R s1 s2.

(**
  Next three lemmas show the two definitions above are strongly related.
*)

    Lemma input_valid_transition_valid
      (l : label)
      (som : state * option message)
      (som' : state * option message)
      (Ht : input_valid_transition l som som')
      : input_valid l som.
    Proof.
      destruct Ht as [Hpv Ht].
      assumption.
    Qed.

    Lemma input_valid_can_transition
      (l : label)
      (som : state * option message)
      (Hv : input_valid l som)
      : forall som', transition l som = som' ->
        input_valid_transition l som som'.
    Proof.
      repeat split; assumption.
    Qed.

    Lemma input_valid_transition_iff
      (l : label)
      (som : state * option message)
      : input_valid l som
      <-> exists (som' : state * option message),
            input_valid_transition l som som'.
    Proof.
      split.
      - eexists.
        apply input_valid_can_transition; [assumption|reflexivity].
      - intros [som' Hivt].
        apply input_valid_transition_valid with som'.
        assumption.
    Qed.

(**

The next couple of lemmas relate the two definitions above with
pre-existing concepts.

 *)
    Lemma input_valid_transition_origin
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s',om'))
      : valid_state_prop s.
    Proof.
      destruct Ht as [[[_om Hp] _] _]. exists _om. assumption.
    Qed.

    Lemma input_valid_transition_destination
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s', om'))
      : valid_state_prop s'.
    Proof.
      exists om'.
      destruct Ht as [[[_om Hs] [[_s Hom] Hv]] Ht].
      apply valid_generated_state_message with s _om _s om l; assumption.
    Qed.

    Lemma input_valid_transition_in
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s', om'))
      : option_valid_message_prop om.
    Proof.
      destruct Ht as [[_ [[_s Hom] _]] _].
      exists _s. assumption.
    Qed.

    Lemma input_valid_transition_outputs_valid_state_message
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s', om'))
        : valid_state_message_prop s' om'.
    Proof.
      destruct Ht as [[[_om Hps] [[_s Hpm] Hv]] Ht].
      apply valid_generated_state_message with s _om _s om l; assumption.
    Qed.

    Lemma input_valid_transition_out
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s', om'))
      : option_valid_message_prop om'.
    Proof.
      apply input_valid_transition_outputs_valid_state_message in Ht.
      exists s'. assumption.
    Qed.

    Lemma input_valid_transition_is_valid
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s', om'))
      : valid l (s, om).
    Proof.
      destruct Ht as [[_ [_ Hv]] _].
      assumption.
    Qed.

    Lemma input_valid_transition_transition
          {l : label}
          {s s' : state}
          {om om' : option message}
          (Ht : input_valid_transition l (s, om) (s', om'))
        :  transition l (s, om) = (s', om').
     Proof.
      destruct Ht as [_ Ht]. assumption.
     Qed.

    Lemma input_valid_state_message_outputs
      (l : label)
      (s : state)
      (om : option message)
      (Hv : input_valid l (s, om))
      s' om'
      (Ht : transition l (s, om) = (s', om'))
      : valid_state_message_prop s' om'.
    Proof.
      destruct Hv as [[_om Hs] [[_s Hom] Hv]].
      apply valid_generated_state_message with s _om _s om l; assumption.
    Qed.

    (** For VLSMs initialized with many initial messages such as
    the [composite_vlsm_constrained_projection] or the [pre_loaded_with_all_messages_vlsm],
    the question of whether a [VLSM] [can_emit] a message <<m>> becomes more
    useful than that whether <<m>> is a [valid_message].
    *)

    Definition option_can_produce
      (s : state)
      (om : option message)
      :=
      exists
      (som : state * option message)
      (l : label),
      input_valid_transition l som (s, om).

    Definition can_produce
      (s : state)
      (m : message)
      := option_can_produce s (Some m).

    (** Of course, if a VLSM [can_emit] <<(s,m)>>, then <<(s,m)>> is valid.
    *)

    Lemma option_can_produce_valid
      (s : state)
      (om : option message)
      (Hm : option_can_produce s om)
      : valid_state_message_prop s om .
    Proof.
      destruct Hm as [(s0, om0) [l [[[_om0 Hs0] [[_s0 Hom0] Hv]] Ht]]].
      apply valid_generated_state_message with s0 _om0 _s0 om0 l; assumption.
    Qed.

    Definition can_produce_valid
      (s : state)
      (m : message)
      (Hm : can_produce s m)
      : valid_state_message_prop s (Some m)
      := option_can_produce_valid s (Some m) Hm.

    Lemma option_can_produce_valid_iff
      (s : state)
      (om : option message)
      : valid_state_message_prop s om <->
        option_can_produce s om \/ initial_state_prop s /\ option_initial_message_prop om.
    Proof.
      split.
      - intros Hm; inversion Hm; subst.
        + right. split; assumption.
        + left.
          exists (s1, om0). exists l0.
          repeat split; [..|assumption|assumption]
          ; eexists; [exact Hps|exact Hpm].
      - intros [Hem | Him].
        + apply option_can_produce_valid. assumption.
        + constructor; apply Him.
    Qed.

    Definition can_produce_valid_iff
      (s : state)
      (m : message)
      : valid_state_message_prop s (Some m) <->
        can_produce s m \/ initial_state_prop s /\ initial_message_prop m
      := option_can_produce_valid_iff s (Some m).

    Definition can_emit
      (m : message)
      :=
      exists
      (som : state * option message)
      (l : label)
      (s : state),
      input_valid_transition l som (s, Some m).

    Lemma can_emit_iff
      (m : message)
      : can_emit m <-> exists s, can_produce s m.
    Proof.
      split.
      - intros [som [l [s Ht]]]. exists s, som, l. assumption.
      - intros [s [som [l Ht]]]. exists som, l, s. assumption.
    Qed.

    (** If a VLSM [can_emit] a message <<m>>, then <<m>> is valid.
    *)

    Lemma emitted_messages_are_valid
      (m : message)
      (Hm : can_emit m)
      : valid_message_prop m .
    Proof.
      apply can_emit_iff in Hm.
      destruct Hm as [s Hm].
      apply can_produce_valid in Hm.
      exists s. assumption.
    Qed.

    (** A characterization of valid messages in terms of [can_emit]
    *)

    Lemma emitted_messages_are_valid_iff
      (m : message)
      : valid_message_prop m <-> initial_message_prop m \/ can_emit m.
    Proof.
      split.
      - intros [s Hm].
        apply can_produce_valid_iff in Hm as [Hgen | [_ Him]].
        + right. apply can_emit_iff. exists s. assumption.
        + left. assumption.
      - intros [Him | Hm].
        + apply initial_message_is_valid. assumption.
        + apply emitted_messages_are_valid. assumption.
    Qed.

(** *** valid state and valid message characterization

The definition and results below show that the mutually-recursive definitions
for [valid_state]s and [valid_message]s can be derived from the
prior definitions.

The results below offers equivalent characterizations for [valid_state]s
and [valid_message]s, similar to their recursive definition.
*)

    Lemma valid_state_prop_iff :
      forall s' : state,
        valid_state_prop s'
        <-> (exists is : initial_state, s' = proj1_sig is)
          \/ exists (l : label) (som : state * option message) (om' : option message),
            input_valid_transition l som (s', om').
    Proof.
      intros; split.
      - intro Hps'. destruct Hps' as [om' Hs].
        inversion Hs; subst.
        * left. exists (exist _ _ Hs0). reflexivity.
        * right. exists l0. exists (s, om). exists om'.
          repeat split; try assumption.
          + exists _om. assumption.
          + exists _s. assumption.
      - intros [[[s His] Heq] | [l [[s om] [om' [[[_om Hps] [[_s Hpm] Hv]] Ht]]]]]; subst.
        + exists None. apply valid_initial_state_message; [assumption | exact I].
        + exists om'. apply valid_generated_state_message with s _om _s om l; assumption.
    Qed.

    (** A specialized induction principle for [valid_state_prop].

        Compared to opening the existential and using [valid_state_message_prop_ind],
        this expresses the inductive assumptions simply in terms of
        [input_valid_transition], rather than than having everything exploded
        as [valid_state_message_prop] assumptions over witnesses <<_s>>
        and <<_om>>, and a spurious inductive assumption <<P _s>>.
     *)
    Lemma valid_state_prop_ind
      (P : state -> Prop)
      (IHinit : forall (s : state) (Hs : initial_state_prop s), P s)
      (IHgen :
        forall (s' : state) (l: label) (om om' : option message) (s : state)
          (Ht : input_valid_transition l (s, om) (s', om')) (Hs : P s),
          P s'
      )
      : forall (s : state) (Hs : valid_state_prop s), P s.
    Proof.
      intros.
      destruct Hs as [om Hs].
      induction Hs.
      - apply IHinit. assumption.
      - apply (IHgen s' l0 om om' s);firstorder.
    Qed.

    (* valid message characterization - similar to the definition in the report. *)

    Lemma valid_message_prop_iff :
      forall m' : message,
        valid_message_prop m'
        <-> (exists im : initial_message, m' = proj1_sig im)
          \/ exists (l : label) (som : state * option message) (s' : state),
            input_valid_transition l som (s', Some m').
    Proof.
      intros; split.
      - intros [s' Hpm'].
        inversion Hpm'; subst.
        + left. exists (exist _ m' Hom). reflexivity.
        + right. exists l0. exists (s, om). exists s'.
          firstorder.
      - intros [[[s His] Heq] | [l [[s om] [s' [[[_om Hps] [[_s Hpm] Hv]] Ht]]]]]; subst.
        + apply initial_message_is_valid. assumption.
        + exists s'.
          apply valid_generated_state_message with s _om _s om l; assumption.
    Qed.

(** ** Trace Properties

Note that it is unnecessary to specify the source state of the transition,
as it is implied by the preceding [transition_item] (or by the <<start>> state,
if such an item doesn't exist).
*)

(**
We will now split our groundwork for defining traces into the finite case and
the infinite case.
*)

(** *** Finite [valid_trace]s

A [finite_valid_trace_from] a [state] <<start>> is a pair <<(start, steps)>> where <<steps>>
is a list of [transition_item]s, and is inductively defined by:
- <<(s, [])>> is a [finite_valid_trace_from] <<s>> if <<s>> is valid
- if there is an [input_valid_transition] <<l (s', iom) (s, oom)>>

  and if <<(s,steps)>> is a [valid_trace_from] <<s>>

  then <<(s', ({| l := l; input := iom; destination := s; output := oom |} :: steps)>>
  is a [finite_valid_trace_from] <<s'>>.

Note that the definition is given such that it extends an existing trace by
adding a transition to its front.
The reason for this choice is to have this definition be similar to the one
for infinite traces, which can only be extended at the front.
*)

    Inductive finite_valid_trace_from : state -> list transition_item -> Prop :=
    | finite_valid_trace_from_empty : forall (s : state)
        (Hs : valid_state_prop s),
        finite_valid_trace_from s []
    | finite_valid_trace_from_extend : forall  (s : state) (tl : list transition_item)
        (Htl : finite_valid_trace_from s tl)
        (s' : state) (iom oom : option message) (l : label)
        (Ht : input_valid_transition l (s', iom) (s, oom)),
        finite_valid_trace_from  s' ({| l := l; input := iom; destination := s; output := oom |} :: tl).

    Definition finite_valid_trace_singleton :
      forall {l : label} {s s': state} {iom oom : option message},
        input_valid_transition l (s, iom) (s', oom) ->
        finite_valid_trace_from  s ({| l := l; input := iom; destination := s'; output := oom |} :: [])
      := fun l s s' iom oom Hptrans =>
           finite_valid_trace_from_extend s' []
               (finite_valid_trace_from_empty s' (input_valid_transition_destination Hptrans))
               _ _ _ _ Hptrans.

(**
To complete our definition of a finite valid trace, we must also guarantee that <<start>> is an
initial state according to the protocol.
*)

    Definition finite_valid_trace (s : state) (ls : list transition_item) : Prop :=
      finite_valid_trace_from s ls /\ initial_state_prop s.

    Opaque finite_valid_trace.

(**
In the remainder of the section we provide various results allowing us to
prove or decompose the above properties in proofs.
*)

    (** This is a bit more useful than the small proof suggests,
        because applying it always leaves just one subgoal.
        The tactical <<split;[constructor;apply initial_state_is_valid|];assumption>>
        only works if the assumption is available, which may require
        an <<assert>> and writing out the full VLSM and state expressions
        as part of the proof script.
     *)
    Lemma finite_valid_trace_empty (s : state):
      vinitial_state_prop X s ->
      finite_valid_trace s [].
    Proof.
      split;[constructor;apply initial_state_is_valid|];assumption.
    Qed.

    Lemma finite_valid_trace_first_valid_transition
          (s : state)
          (tr : list transition_item)
          (te : transition_item)
          (Htr : finite_valid_trace_from s (te :: tr))
      : input_valid_transition (l te) (s, input te) (destination te, output te).
    Proof.
      inversion Htr. assumption.
    Qed.

    Lemma finite_valid_trace_first_pstate
      (s : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from s tr)
      : valid_state_prop s.
    Proof.
      inversion Htr; subst; [assumption|].
      apply Ht.
    Qed.

    Lemma finite_valid_trace_tail
          (s : state)
          (tr : list transition_item)
          (te : transition_item)
          (Htr : finite_valid_trace_from s (te :: tr))
      : finite_valid_trace_from (destination te) tr.
    Proof.
      inversion Htr. assumption.
    Qed.

    Lemma finite_valid_trace_last_pstate
      (s : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from s tr)
      : valid_state_prop (finite_trace_last s tr).
    Proof.
      generalize dependent s.
      induction tr; intros.
      - simpl. apply finite_valid_trace_first_pstate with []. assumption.
      - apply finite_valid_trace_tail in Htr.
        apply IHtr in Htr.
        replace
          (finite_trace_last s (a :: tr))
          with (finite_trace_last (destination a) tr)
        ;[assumption|].
        unfold finite_trace_last.
        rewrite map_cons.
        rewrite unroll_last.
        reflexivity.
    Qed.

    Lemma input_valid_transition_to
          (s : state)
          (tr : list transition_item)
          (tr1 tr2 : list transition_item)
          (te : transition_item)
          (Htr : finite_valid_trace_from s tr)
          (Heq : tr = tr1 ++ [te] ++ tr2)
          (lst1 := finite_trace_last s tr1)
      : input_valid_transition (l te) (lst1, input te) (destination te, output te).
    Proof.
      generalize dependent s. generalize dependent tr.
      induction tr1.
      - intros tr Heq s Htr. simpl in Heq; subst. inversion Htr; subst. assumption.
      - specialize (IHtr1 (tr1 ++ [te] ++ tr2) eq_refl).
        intros tr Heq is Htr; subst. inversion Htr; subst.
        rewrite finite_trace_last_cons.
        apply IHtr1. assumption.
    Qed.

    Lemma finite_valid_trace_consecutive_valid_transition
          (s : state)
          (tr : list transition_item)
          (tr1 tr2 : list transition_item)
          (te1 te2 : transition_item)
          (Htr : finite_valid_trace_from s tr)
          (Heq : tr = tr1 ++ [te1; te2] ++ tr2)
      : input_valid_transition (l te2) (destination te1, input te2) (destination te2, output te2).
    Proof.
      change ([te1; te2] ++ tr2) with ([te1] ++ [te2] ++ tr2) in Heq.
      rewrite app_assoc in Heq.
      specialize (input_valid_transition_to s tr (tr1 ++ [te1]) tr2 te2 Htr Heq)
        as Ht.
      rewrite finite_trace_last_is_last in Ht. assumption.
    Qed.


    Lemma valid_trace_output_is_valid
      (is : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from is tr)
      (m : message)
      (Houtput : trace_has_message (field_selector output) m tr)
      : valid_message_prop m.
    Proof.
      revert is Htr.
      induction Houtput as [item tr' Hm| item tr'];intros;inversion Htr; subst.
      - simpl in Hm.
        subst.
        apply input_valid_transition_out in Ht.
        assumption.
      - apply (IHHoutput s).
        assumption.
    Qed.

    Lemma valid_trace_input_is_valid
      (is : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from is tr)
      (m : message)
      (Hinput : trace_has_message (field_selector input) m tr)
      : valid_message_prop m.
    Proof.
      revert is Htr.
      induction Hinput as [item tr' Hm| item tr'];intros
      ;inversion Htr as [|s _tr'  Htr' _is iom oom l Ht ];subst.
      - simpl in Hm.
        subst.
        apply input_valid_transition_in in Ht.
        assumption.
      - apply (IHHinput s).
        assumption.
    Qed.

    Lemma valid_trace_observed_is_valid
      (is : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from is tr)
      (m : message)
      (Hobserved : trace_has_message item_sends_or_receives m tr)
      : valid_message_prop m.
    Proof.
      apply trace_has_message_observed_iff in Hobserved as [Hm |Hm]
      ; revert Htr m Hm; [apply valid_trace_input_is_valid | apply valid_trace_output_is_valid].
    Qed.

    Lemma first_transition_valid
      (s : state)
      (te : transition_item)
      : finite_valid_trace_from s [te] <-> input_valid_transition (l te) (s, input te) (destination te, output te).

    Proof.
      split.
      - intro Htr.
        inversion Htr.
        assumption.
      - destruct te. simpl. intro Ht.
        apply input_valid_transition_destination in Ht as Hdestination0.
        constructor; [|assumption]. constructor. assumption.
    Qed.

    Lemma extend_right_finite_trace_from
      (s1 : state)
      (ts : list transition_item)
      (Ht12 : finite_valid_trace_from s1 ts)
      (l3 : label)
      (s2 := finite_trace_last s1 ts)
      (iom3 : option message)
      (s3 : state)
      (oom3 : option message)
      (Hv23 : input_valid_transition l3 (s2, iom3) (s3, oom3))
      : finite_valid_trace_from s1 (ts ++ [{| l := l3; destination := s3; input := iom3; output := oom3 |}]).
    Proof.
      induction Ht12.
      - simpl. apply finite_valid_trace_singleton;assumption.
      - rewrite <- app_comm_cons.
        apply finite_valid_trace_from_extend; try assumption.
        simpl in IHHt12. apply IHHt12.
        unfold s2 in *; clear s2.
        rewrite finite_trace_last_cons in Hv23.
        assumption.
    Qed.

(**
We can now prove several general properties of [finite_valid_trace]s. For example,
the following lemma states that given two such traces, such that the latter's starting state
is equal to the former's last state, it is possible to _concatenate_ them into a single
[finite_valid_trace].
*)

    Lemma finite_valid_trace_from_app_iff (s : state) (ls ls' : list transition_item) (s' := finite_trace_last s ls)
      : finite_valid_trace_from s ls /\ finite_valid_trace_from s' ls'
        <->
        finite_valid_trace_from s (ls ++ ls').
    Proof.
      subst s'.
      revert s.
      induction ls;intro s.
      - rewrite finite_trace_last_nil. simpl.
        intuition (eauto using finite_valid_trace_first_pstate, finite_valid_trace_from_empty).
      - rewrite finite_trace_last_cons. simpl.
        specialize (IHls (destination a)).
        split.
        + intros [Hal Hl'].
          inversion Hal; subst; simpl in *.
          constructor;[apply IHls;split|];assumption.
        + inversion 1;subst; simpl in *.
          apply IHls in Htl as [Hl Hl'].
          split;[constructor|];assumption.
    Qed.

    Lemma finite_valid_trace_from_rev_ind
      (P : state -> list transition_item -> Prop)
      (Hempty: forall s,
        valid_state_prop s -> P s nil)
      (Hextend : forall s tr,
        finite_valid_trace_from s tr ->
        P s tr ->
        forall sf iom oom l
        (Hx: input_valid_transition l (finite_trace_last s tr,iom) (sf,oom)),
        let x:= {|l:=l; input:=iom; destination:=sf; output:=oom|} in
        P s (tr++[x])):
      forall s tr,
        finite_valid_trace_from s tr ->
        P s tr.
    Proof.
      induction tr using rev_ind; intro Htr.
      - inversion Htr. apply Hempty. congruence.
      - apply finite_valid_trace_from_app_iff in Htr.
        destruct Htr as [Htr Hx].
        destruct x; apply (Hextend _ _ Htr (IHtr Htr)).
        inversion Hx; congruence.
    Qed.

    Lemma finite_valid_trace_rev_ind
      (P : state -> list transition_item -> Prop)
      (Hempty: forall si,
        initial_state_prop si -> P si nil)
      (Hextend : forall si tr,
        finite_valid_trace si tr ->
        P si tr ->
        forall sf iom oom l
        (Hx: input_valid_transition l (finite_trace_last si tr,iom) (sf,oom)),
        let x:= {|l:=l; input:=iom; destination:=sf; output:=oom|} in
        P si (tr++[x])):
      forall si tr,
        finite_valid_trace si tr ->
        P si tr.
    Proof.
      intros si tr [Htr Hinit].
      induction Htr using finite_valid_trace_from_rev_ind.
      - apply Hempty;auto.
      - apply Hextend;[split|..];auto.
    Qed.

(** Several other lemmas in this vein are necessary for proving results regarding
traces.
*)

    Lemma finite_valid_trace_from_prefix
      (s : state)
      (ls : list transition_item)
      (Htr : finite_valid_trace_from s ls)
      (n : nat)
      : finite_valid_trace_from s (list_prefix ls n).
    Proof.
      specialize (list_prefix_suffix ls n); intro Hdecompose.
      rewrite <- Hdecompose in Htr.
      apply finite_valid_trace_from_app_iff in Htr.
      destruct Htr as [Hpr _].
      assumption.
    Qed.

    Lemma finite_valid_trace_from_suffix
      (s : state)
      (ls : list transition_item)
      (Htr : finite_valid_trace_from s ls)
      (n : nat)
      (nth : state)
      (Hnth : finite_trace_nth s ls n = Some nth)
      : finite_valid_trace_from nth (list_suffix ls n).
    Proof.
      rewrite <- (list_prefix_suffix ls n) in Htr.
      apply finite_valid_trace_from_app_iff in Htr.
      destruct Htr as [_ Htr].
      replace (finite_trace_last s (list_prefix ls n)) with nth in Htr;[assumption|].
      {
        destruct n.
        - rewrite finite_trace_nth_first in Hnth. injection Hnth as ->.
          destruct ls;reflexivity.
        - unfold finite_trace_last.
          rewrite list_prefix_map.
          apply list_prefix_nth_last.
          assumption.
      }
    Qed.

    Lemma finite_valid_trace_from_segment
      (s : state)
      (ls : list transition_item)
      (Htr : finite_valid_trace_from s ls)
      (n1 n2 : nat)
      (Hle : n1 <= n2)
      (n1th : state)
      (Hnth : finite_trace_nth s ls n1 = Some n1th)
      : finite_valid_trace_from n1th (list_segment ls n1 n2).
    Proof.
      apply finite_valid_trace_from_suffix with s.
      - apply finite_valid_trace_from_prefix. assumption.
      - destruct n1;[assumption|].
        unfold finite_trace_nth in Hnth |- *.
        simpl in Hnth |- *.
        rewrite list_prefix_map.
        rewrite list_prefix_nth;assumption.
    Qed.

    (* begin hide *)

    Lemma can_produce_from_valid_trace si tr
      (Htr: finite_valid_trace_from si tr)
      : forall item, item ∈ tr ->
        option_can_produce (destination item) (output item).
    Proof.
      intros item Hitem.
      apply elem_of_list_split in Hitem as (l1 & l2 & Heq).
      eexists _,_.
      eapply input_valid_transition_to; [eassumption|].
      simpl. eassumption.
    Qed.

    Lemma can_emit_from_valid_trace
      (si : state)
      (m : message)
      (tr : list transition_item)
      (Htr: finite_valid_trace si tr)
      (Hm : trace_has_message (field_selector output) m tr) :
      can_emit m.
    Proof.
      apply can_emit_iff.
      revert Hm.
      setoid_rewrite Exists_exists.
      intros [item [Hitem Houtput]].
      exists (destination item).
      unfold can_produce.
      replace (Some m) with (output item) by assumption.
      eapply can_produce_from_valid_trace; [apply Htr|assumption].
    Qed.

    (* End Hide *)

(**
** Finite [valid_trace]s with a final state
*)

(**
It is often necessary to refer to know ending state of a [finite_valid_trace_from].
This is either the [destination] of the [last] [transition_item] in the trace, or
the starting state.
To avoid repeating reasoning about [last], we define variants of
[finite_valid_trace_from] and [finite_valid_trace]
that include the final state, and give appropriate induction principles.
 *)

(** The final state of a finite portion of a valid trace.
    This is defined over [finite_valid_trace_from] because
    an initial state is necessary in case <<tr>> is empty,
    and this allows the definition to have only one non-implicit
    parameter.
 *)

    Inductive finite_valid_trace_from_to : state -> state -> list transition_item -> Prop :=
    | finite_valid_trace_from_to_empty : forall (s : state)
        (Hs : valid_state_prop s),
        finite_valid_trace_from_to s s []
    | finite_valid_trace_from_to_extend : forall  (s f : state) (tl : list transition_item)
        (Htl : finite_valid_trace_from_to s f tl)
        (s' : state) (iom oom : option message) (l : label)
        (Ht : input_valid_transition l (s', iom) (s, oom)),
        finite_valid_trace_from_to s' f ({| l := l; input := iom; destination := s; output := oom |} :: tl).

    Lemma finite_valid_trace_from_to_singleton s s' iom oom l
        : input_valid_transition l (s, iom) (s', oom) ->
          finite_valid_trace_from_to s s' [{| l := l; input := iom; destination := s'; output := oom |}].
    Proof.
      intro Ht.
      constructor;[|assumption].
      constructor.
      apply input_valid_transition_destination in Ht.
      assumption.
    Qed.

    Lemma finite_valid_trace_from_to_forget_last
          s f tr : finite_valid_trace_from_to s f tr -> finite_valid_trace_from s tr.
    Proof.
      induction 1;constructor;auto.
    Qed.

    Lemma finite_valid_trace_from_to_last
          s f tr : finite_valid_trace_from_to s f tr -> finite_trace_last s tr = f.
    Proof.
      induction 1.
      - apply finite_trace_last_nil.
      - rewrite finite_trace_last_cons; assumption.
    Qed.


    Lemma finite_valid_trace_from_add_last
          s f tr :
      finite_valid_trace_from s tr ->
      finite_trace_last s tr = f ->
      finite_valid_trace_from_to s f tr.
    Proof.
      intro Hfrom.
      induction Hfrom.
      - rewrite finite_trace_last_nil. intros <-.
        constructor. assumption.
      - rewrite finite_trace_last_cons. simpl. intro.
        constructor;auto.
    Qed.

    Lemma finite_valid_trace_from_to_first_pstate
          s f tr : finite_valid_trace_from_to s f tr -> valid_state_prop s.
    Proof.
      intro Htr.
      apply finite_valid_trace_from_to_forget_last in Htr.
      apply finite_valid_trace_first_pstate in Htr.
      assumption.
    Qed.

    Lemma finite_valid_trace_from_to_last_pstate
          s f tr : finite_valid_trace_from_to s f tr -> valid_state_prop f.
    Proof.
      intro Htr.
      rewrite <- (finite_valid_trace_from_to_last _ _ _ Htr).
      apply finite_valid_trace_last_pstate.
      apply finite_valid_trace_from_to_forget_last in Htr.
      assumption.
    Qed.

    Lemma finite_valid_trace_from_to_app
      (m s f: state) (ls ls' : list transition_item)
      : finite_valid_trace_from_to s m ls
        -> finite_valid_trace_from_to m f ls'
        -> finite_valid_trace_from_to s f (ls ++ ls').
    Proof.
      intros Hl Hl';induction Hl;simpl.
      - trivial.
      - constructor;auto.
    Qed.

    Lemma finite_valid_trace_from_to_app_split
      (s f: state) (ls ls' : list transition_item)
      : finite_valid_trace_from_to s f (ls ++ ls') ->
        let m := finite_trace_last s ls in
        finite_valid_trace_from_to s m ls
        /\ finite_valid_trace_from_to m f ls'.
    Proof.
      revert s;induction ls;intros s;simpl.
      - rewrite finite_trace_last_nil.
        intro Htr. split;[|assumption].
        apply finite_valid_trace_from_to_first_pstate in Htr.
        constructor;assumption.
      - rewrite finite_trace_last_cons.
        inversion 1; subst; simpl in *.
        apply IHls in Htl as [].
        auto using finite_valid_trace_from_to_extend.
    Qed.

    Definition finite_valid_trace_init_to si sf tr : Prop
      := finite_valid_trace_from_to si sf tr
          /\ initial_state_prop si.

    Lemma finite_valid_trace_init_add_last si sf tr:
      finite_valid_trace si tr ->
      finite_trace_last si tr = sf ->
      finite_valid_trace_init_to si sf tr.
    Proof.
      intros [Htr Hinit] Hf.
      split;eauto using finite_valid_trace_from_add_last.
    Qed.

    Lemma finite_valid_trace_init_to_forget_last si sf tr:
      finite_valid_trace_init_to si sf tr ->
      finite_valid_trace si tr.
    Proof.
      intros [Hinit Htr].
      split;eauto using finite_valid_trace_from_to_forget_last.
    Qed.

    Lemma finite_valid_trace_init_to_last si sf tr:
      finite_valid_trace_init_to si sf tr ->
      finite_trace_last si tr = sf.
    Proof.
      intros [Htr _].
      eauto using finite_valid_trace_from_to_last.
    Qed.

    Lemma extend_right_finite_trace_from_to
      (s1 s2 : state)
      (ts : list transition_item)
      (Ht12 : finite_valid_trace_from_to s1 s2 ts)
      (l3 : label)
      (iom3 : option message)
      (s3 : state)
      (oom3 : option message)
      (Hv23 : input_valid_transition l3 (s2, iom3) (s3, oom3))
      : finite_valid_trace_from_to s1 s3 (ts ++ [{| l := l3; destination := s3; input := iom3; output := oom3 |}]).
    Proof.
      induction Ht12.
      - simpl. apply finite_valid_trace_from_to_singleton;assumption.
      - rewrite <- app_comm_cons.
        apply finite_valid_trace_from_to_extend; auto.
    Qed.

    Lemma finite_valid_trace_from_to_rev_ind
      (P : state -> state -> list transition_item -> Prop)
      (Hempty: forall si
        (Hsi : valid_state_prop si),
        P si si nil)
      (Hextend : forall si s tr
        (IHtr : P si s tr)
        (Htr : finite_valid_trace_from_to si s tr)
        sf iom oom l
        (Ht : input_valid_transition l (s,iom) (sf,oom)),
        P si sf (tr++[{|l:=l; input:=iom; destination:=sf; output:=oom|}])):
      forall si sf tr,
        finite_valid_trace_from_to si sf tr ->
        P si sf tr.
    Proof.
      intros si sf tr Htr.
      revert sf Htr.
      induction tr using rev_ind;
      intros sf Htr.
      - inversion Htr;subst. apply Hempty;assumption.
      - apply finite_valid_trace_from_to_app_split in Htr.
        destruct Htr as [Htr Hstep].
        inversion Hstep;subst.
        inversion Htl;subst.
        revert Ht.
        apply Hextend; [|assumption].
        apply IHtr.
        assumption.
    Qed.

    Lemma finite_valid_trace_init_to_rev_ind
      (P : state -> state -> list transition_item -> Prop)
      (Hempty: forall si
        (Hsi : initial_state_prop si),
        P si si nil)
      (Hextend : forall si s tr
        (IHtr : P si s tr)
        (Htr : finite_valid_trace_init_to si s tr)
        sf iom oom l
        (Ht : input_valid_transition l (s,iom) (sf,oom)),
        P si sf (tr++[{|l:=l; input:=iom; destination:=sf; output:=oom|}])):
      forall si sf tr,
        finite_valid_trace_init_to si sf tr ->
        P si sf tr.
    Proof.
      intros si sf tr Htr.
      destruct Htr as [Htr Hinit].
      induction Htr using finite_valid_trace_from_to_rev_ind.
      - apply Hempty. assumption.
      - apply Hextend with s.
        + apply IHHtr. assumption.
        + split; assumption.
        + assumption.
    Qed.

(** An inductive valid trace property which also identifies the final message.

As shown by the [finite_valid_trace_init_to_emit_valid_state_message]  and
[finite_valid_trace_init_to_emit_valid_state_message_rev] lemmas below, this definition
is the trace-equivalent of the [valid_state_message_prop]erty.

This inductive property is reflecting that fact that a that <<valid_state_message_prop (s,om)>>
holds only if <<s>> and <<om>> are the final state and output of an initial valid
trace, or a pair of an initial state and option-initial message.
It follows the inductive structure of <<valid_state_message_prop>>, but augments every node of
the tree with such an exhibiting trace.

Its main benefit is that when performing induction over it, one can also use the
induction hypothesis for the (trace generating the) message being received.

Although this definition could be used directly, we prefer to use it to derive
a stronger induction principle ([finite_valid_trace_init_to_rev_strong_ind])
over [finite_valid_trace_init_to] traces.
*)
    Inductive finite_valid_trace_init_to_emit : state -> state -> option message -> list transition_item -> Prop :=
    | finite_valid_trace_init_to_emit_empty : forall (is : state) (om : option message)
        (His : initial_state_prop is)
        (Him : option_initial_message_prop om),
        finite_valid_trace_init_to_emit is is om []
    | finite_valid_trace_init_to_emit_extend
        : forall
          (is s : state) (_om : option message) (tl : list transition_item)
          (Hs : finite_valid_trace_init_to_emit is s _om tl)
          (iom_is iom_s : state) (iom : option message) (iom_tl : list transition_item)
          (Hiom : finite_valid_trace_init_to_emit iom_is iom_s iom iom_tl)
          (l : label)
          (Hv : valid l (s, iom))
          (s' : state) (oom : option message)
          (Ht : transition l (s, iom) = (s', oom)),
          finite_valid_trace_init_to_emit is s' oom (tl ++ [{| l := l; input := iom; destination := s'; output := oom |}]).

    Lemma finite_valid_trace_init_to_emit_initial_state
      (is f : state) (om : option message) (tl : list transition_item)
      (Htl : finite_valid_trace_init_to_emit is f om tl)
      : initial_state_prop is.
    Proof.
      induction Htl; assumption.
    Qed.

(** A property characterizing the "emit" message of [finite_valid_trace_init_to_emit].

There are two cases: (1) either the trace is empty, and then we require
the message to be initial; or (2) the trace is not empty, and the message
is the output of the last transition.
*)
    Definition empty_initial_message_or_final_output (tl : list transition_item) (om : option message) : Prop.
    Proof.
      destruct (has_last_or_null tl) as [[_ [item _]] | _].
      - exact (output item  = om).
      - exact (option_initial_message_prop om).
    Defined.

    Lemma finite_valid_trace_init_to_emit_output
      (s f : state) (om : option message) (tl : list transition_item)
      (Htl : finite_valid_trace_init_to_emit s f om tl)
      : empty_initial_message_or_final_output tl om.
    Proof.
      unfold empty_initial_message_or_final_output.
      destruct_list_last tl tl' item Heqtl.
      - inversion Htl; [assumption|].
        destruct tl0; simpl in *; congruence.
      - rewrite <- Heqtl in Htl.
        inversion Htl; [destruct tl'; simpl in *; congruence|].
        revert Heqtl; subst; intro Heqtl.
        apply app_inj_tail, proj2 in Heqtl. subst. reflexivity.
    Qed.

    Lemma finite_valid_trace_init_to_emit_valid_state_message
      (s f : state) (om : option message) (tl : list transition_item)
      (Htl : finite_valid_trace_init_to_emit s f om tl)
      : valid_state_message_prop f om.
    Proof.
      induction Htl.
      - apply valid_initial_state_message; assumption.
      - apply valid_generated_state_message with s _om iom_s iom l0; assumption.
    Qed.

    Lemma finite_valid_trace_init_to_emit_valid_state_message_rev
      f om
      (Hp : valid_state_message_prop f om)
      : exists (s : state) (tl : list transition_item),
        finite_valid_trace_init_to_emit s f om tl.
    Proof.
      induction Hp.
      - exists s, []. constructor; assumption.
      - destruct IHHp1 as [is [tl Hs]].
        destruct IHHp2 as [om_is [om_tl Hom]].
        eexists; eexists.
        apply
          (finite_valid_trace_init_to_emit_extend _ _ _ _ Hs _ _ _ _ Hom _ Hv _ _ Ht).
    Qed.

    Lemma finite_valid_trace_init_to_emit_forget_emit
      (s f : state) (_om : option message) (tl : list transition_item)
      (Htl : finite_valid_trace_init_to_emit s f _om tl)
      : finite_valid_trace_init_to s f tl.
    Proof.
      apply finite_valid_trace_init_to_emit_initial_state in Htl as Hinit.
      split; [|assumption].
      clear Hinit.
      induction Htl.
      - constructor. apply initial_state_is_valid. assumption.
      - apply finite_valid_trace_from_to_app with s; [assumption|].
        apply finite_valid_trace_from_to_singleton.
        apply finite_valid_trace_init_to_emit_valid_state_message in Htl1.
        apply finite_valid_trace_init_to_emit_valid_state_message in Htl2.
        repeat split; [..|assumption|assumption]; eexists; [exact Htl1 | exact Htl2].
    Qed.

    Lemma finite_valid_trace_init_to_add_emit
      (s f : state) (tl : list transition_item)
      (Htl : finite_valid_trace_init_to s f tl)
      : finite_valid_trace_init_to_emit s f (finite_trace_last_output tl) tl.
    Proof.
      induction Htl using finite_valid_trace_init_to_rev_ind.
      - constructor; [assumption | exact I].
      - rewrite finite_trace_last_output_is_last. simpl.
        destruct Ht as [[_ [[_s Hiom] Hv]] Ht].
        specialize (finite_valid_trace_init_to_emit_valid_state_message_rev _ _ Hiom) as [iom_s [iom_tr Hiom_tr]].
        apply (finite_valid_trace_init_to_emit_extend _ _ _ _ IHHtl _ _ _ _ Hiom_tr _ Hv _ _ Ht).
    Qed.

(** Inspired by [finite_valid_trace_init_to_add_emit], we can derive
an induction principle for [finite_valid_trace_init_to] stronger than
[finite_valid_trace_init_to_rev_ind], which allows the induction hypothesis
to be used for the trace generating the message received in the last transition.
*)
    Lemma finite_valid_trace_init_to_rev_strong_ind
      (P : state -> state -> list transition_item -> Prop)
      (Hempty: forall is
        (His : initial_state_prop is),
        P is is nil)
      (Hextend : forall is s tr
        (IHs : P is s tr)
        (Hs : finite_valid_trace_init_to is s tr)
        iom iom_si iom_s iom_tr
        (Heqiom : empty_initial_message_or_final_output iom_tr iom)
        (IHiom : P iom_si iom_s iom_tr)
        (Hiom : finite_valid_trace_init_to iom_si iom_s iom_tr)
        sf oom l
        (Ht : input_valid_transition l (s,iom) (sf,oom)),
        P is sf (tr++[{|l:=l; input:=iom; destination:=sf; output:=oom|}]))
      : forall si sf tr,
        finite_valid_trace_init_to si sf tr ->
        P si sf tr.
    Proof.
      intros is sf tr Htr.
      apply finite_valid_trace_init_to_add_emit in Htr.
      remember (finite_trace_last_output tr) as om. clear Heqom.
      induction Htr.
      - apply Hempty. assumption.
      - assert (Hivt : input_valid_transition l0 (s, iom) (s', oom)).
        { apply finite_valid_trace_init_to_emit_valid_state_message in Htr1.
          apply finite_valid_trace_init_to_emit_valid_state_message in Htr2.
          repeat split; [..|assumption|assumption]; eexists; [exact Htr1 | exact Htr2].
        }
        apply finite_valid_trace_init_to_emit_output in Htr2 as Houtput.
        apply finite_valid_trace_init_to_emit_forget_emit in Htr1.
        apply finite_valid_trace_init_to_emit_forget_emit in Htr2.
        apply (Hextend _ _ _ IHHtr1 Htr1 _ _ _ _ Houtput IHHtr2 Htr2 _ _ _ Hivt).
    Qed.

(** *** Infinite [protcol_trace]s *)

(** We now define [infinite_valid_trace]s. The definitions
resemble their finite counterparts, adapted to the technical
necessities of defining infinite objects. Notably, <<steps>> is
stored as a stream, as opposed to a list.
*)

    CoInductive infinite_valid_trace_from :
      state -> Stream transition_item -> Prop :=
    | infinite_valid_trace_from_extend : forall  (s : state) (tl : Stream transition_item)
        (Htl : infinite_valid_trace_from s tl)
        (s' : state) (iom oom : option message) (l : label)
        (Ht : input_valid_transition l (s', iom) (s, oom)),
        infinite_valid_trace_from  s' (Cons {| l := l; input := iom; destination := s; output := oom |}  tl).

    Definition infinite_valid_trace (s : state) (st : Stream transition_item)
      := infinite_valid_trace_from s st /\ initial_state_prop s.

(**
As for the finite case, the following lemmas help decompose teh above
definitions, mostly reducing them to properties about their finite segments.
*)
    Lemma infinite_valid_trace_consecutive_valid_transition
          (is : state)
          (tr tr2 : Stream transition_item)
          (tr1 : list transition_item)
          (te1 te2 : transition_item)
          (Htr : infinite_valid_trace_from is tr)
          (Heq : tr = stream_app (tr1 ++ [te1; te2]) tr2)
      : input_valid_transition (l te2) (destination te1, input te2) (destination te2, output te2).
    Proof.
      generalize dependent is. generalize dependent tr.
      induction tr1.
      - intros tr Heq is Htr. simpl in Heq; subst. inversion Htr; subst. inversion Htl; subst. assumption.
      - specialize (IHtr1 (stream_app (tr1 ++ [te1; te2]) tr2) eq_refl).
        intros tr Heq is Htr; subst. inversion Htr; subst.
        specialize (IHtr1 s Htl). assumption.
    Qed.

    Lemma infinite_valid_trace_from_app_iff
      (s : state)
      (ls : list transition_item)
      (ls' : Stream transition_item)
      (s' := finite_trace_last s ls)
      : finite_valid_trace_from s ls /\ infinite_valid_trace_from s' ls'
        <->
        infinite_valid_trace_from s (stream_app ls ls').
    Proof.
      intros. generalize dependent ls'. generalize dependent s.
      induction ls; intros; split.
      - destruct 1. assumption.
      - simpl; intros Hls'; split; try assumption. constructor. inversion Hls'; try assumption.
        apply (input_valid_transition_origin Ht).
      - simpl. intros [Htr Htr'].
        destruct a. apply infinite_valid_trace_from_extend.
        + apply IHls. inversion Htr. split. apply Htl.
          unfold s' in Htr'.
          rewrite finite_trace_last_cons in Htr'.
          assumption.
        + inversion Htr. apply Ht.
       - inversion 1. subst. specialize (IHls s1). simpl in IHls. specialize (IHls ls'). apply IHls in Htl.
         destruct Htl. split.
         + constructor; assumption.
         + unfold s'. rewrite finite_trace_last_cons. assumption.
    Qed.

    Lemma infinite_valid_trace_from_prefix
      (s : state)
      (ls : Stream transition_item)
      (Htr : infinite_valid_trace_from s ls)
      (n : nat)
      : finite_valid_trace_from s (stream_prefix ls n).
    Proof.
      specialize (stream_prefix_suffix ls n); intro Hdecompose.
      rewrite <- Hdecompose in Htr.
      apply infinite_valid_trace_from_app_iff in Htr.
      destruct Htr as [Hpr _].
      assumption.
    Qed.

    Lemma infinite_valid_trace_from_prefix_rev
      (s : state)
      (ls : Stream transition_item)
      (Hpref: forall n : nat, finite_valid_trace_from s (stream_prefix ls n))
      : infinite_valid_trace_from s ls.
    Proof.
      revert s ls Hpref.
      cofix Hls.
      intros s (a, ls) Hpref.
      assert (Hpref0 := Hpref 1).
      inversion Hpref0; subst.
      constructor; try assumption.
      apply Hls.
      intro n.
      specialize (Hpref (S n)).
      simpl in Hpref.
      inversion Hpref; subst.
      assumption.
    Qed.

    Lemma infinite_valid_trace_from_EqSt :
      forall s tl1 tl2, EqSt tl1 tl2 -> infinite_valid_trace_from s tl1 -> infinite_valid_trace_from s tl2.
    Proof.
      intros s tl1 tl2 Heq Htl1.
      apply infinite_valid_trace_from_prefix_rev.
      intro n.
      apply stream_prefix_EqSt with (n0 := n) in Heq.
      apply infinite_valid_trace_from_prefix with (n := n) in Htl1.
      rewrite <- Heq. assumption.
    Qed.

    Lemma infinite_valid_trace_from_segment
      (s : state)
      (ls : Stream transition_item)
      (Htr : infinite_valid_trace_from s ls)
      (n1 n2 : nat)
      (Hle : n1 <= n2)
      (n1th := Str_nth n1 (Cons s (Streams.map destination ls)))
      : finite_valid_trace_from n1th (stream_segment ls n1 n2).
    Proof.
      apply finite_valid_trace_from_suffix with s.
      - apply infinite_valid_trace_from_prefix. assumption.
      - destruct n1; try reflexivity.
        unfold n1th. clear n1th.
        unfold finite_trace_nth.
        simpl.
        rewrite stream_prefix_map.
        rewrite stream_prefix_nth; try assumption.
        reflexivity.
    Qed.

(** *** valid traces

Finally, we define [Trace] as a sum-type of its finite/infinite variants.
It inherits some previously introduced definitions, culminating with the
[valid_trace].
*)

    Definition valid_trace_from_prop (tr : Trace) : Prop :=
      match tr with
      | Finite s ls => finite_valid_trace_from s ls
      | Infinite s sm => infinite_valid_trace_from s sm
      end.

    Definition valid_trace_prop (tr : Trace) : Prop :=
      match tr with
      | Finite s ls => finite_valid_trace s ls
      | Infinite s sm => infinite_valid_trace s sm
      end.

    Definition valid_trace : Type :=
      { tr : Trace | valid_trace_prop tr}.

    Lemma valid_trace_from
      (tr : Trace)
      (Htr : valid_trace_prop tr)
      : valid_trace_from_prop tr.
    Proof.
      destruct tr; simpl; destruct Htr as [Htr Hinit]; assumption.
    Qed.

    Lemma valid_trace_initial
      (tr : Trace)
      (Htr : valid_trace_prop tr)
      : initial_state_prop (trace_first tr).
    Proof.
      destruct tr; simpl; destruct Htr as [Htr Hinit]; assumption.
    Qed.

    Lemma valid_trace_from_iff
      (tr : Trace)
      : valid_trace_prop tr
      <-> valid_trace_from_prop tr /\ initial_state_prop (trace_first tr).
    Proof.
      split.
      - intro Htr; split.
        + apply valid_trace_from; assumption.
        + apply valid_trace_initial; assumption.
      - destruct tr; simpl; intros [Htr Hinit]; split; assumption.
    Qed.

(** Having defined [valid_trace]s, we now connect them to valid states
and messages, in the following sense: for each state-message pair (<<s>>, <<m>>)
that has the [valid_state_message_prop]erty, there exists a [valid_trace] which ends
in <<s>> by outputting <<m>> *)

    Lemma valid_state_message_has_trace
          (s : state)
          (om : option message)
          (Hp : valid_state_message_prop s om)
      : initial_state_prop s /\ option_initial_message_prop om
      \/ exists (is : state) (tr : list transition_item),
            finite_valid_trace_init_to is s tr
            /\ finite_trace_last_output tr = om.
    Proof.
      apply finite_valid_trace_init_to_emit_valid_state_message_rev in Hp as [is [tr Htr]].
      apply finite_valid_trace_init_to_emit_output in Htr as Houtput.
      unfold empty_initial_message_or_final_output in Houtput.
      destruct_list_last tr tr' item Heqtr.
      - left. split; [|assumption]. inversion Htr; [assumption|].
        destruct tl; simpl in *; congruence.
      - right. apply finite_valid_trace_init_to_emit_forget_emit in Htr.
        eexists _,_. split; [exact Htr|].
        rewrite finite_trace_last_output_is_last. assumption.
    Qed.

    (** Giving a trace for [valid_state_prop] can be stated more
        simply than [valid_state_message_has_trace], because we don't need a
        disjunction because we are not making claims about [output]
        messages.
     *)
    Lemma valid_state_has_trace
          (s : state)
          (Hp : valid_state_prop s):
      exists (is : state) (tr : list transition_item),
        finite_valid_trace_init_to is s tr.
    Proof using.
      destruct Hp as [_om Hp].
      apply valid_state_message_has_trace in Hp.
      destruct Hp as [[Hinit _]|Htrace].
      + exists s, [].
        split;[|assumption].
        constructor.
        apply initial_state_is_valid.
        assumption.
      + destruct Htrace as [is [tr [Htr _]]].
        exists is, tr.
        assumption.
    Qed.

    (** For any input valid transition there exists a valid trace ending in it. *)
    Lemma exists_right_finite_trace_from
      l s1 iom s2 oom
      (Ht : input_valid_transition l (s1, iom) (s2, oom))
      : exists s0 ts, finite_valid_trace_init_to s0 s2 (ts ++ [{| l := l; destination := s2; input := iom; output := oom |}])
        /\ finite_trace_last s0 ts = s1.
    Proof.
      apply input_valid_transition_origin in Ht as Hs1.
      apply valid_state_has_trace in Hs1.
      destruct Hs1 as [s0 [ts Hts]].
      exists s0, ts.
      destruct Hts as [Hts Hinit].
      repeat split; [|assumption|revert Hts; apply finite_valid_trace_from_to_last].
      revert Ht.
      apply extend_right_finite_trace_from_to.
      assumption.
    Qed.

    Lemma can_emit_has_trace m :
      can_emit m ->
      exists is tr item,
      finite_valid_trace is (tr ++ [item]) /\
      output item = Some m.
    Proof.
      intros [(s, im) [l [s' Hm]]].
      apply exists_right_finite_trace_from in Hm as [is [tr [Htr _]]].
      apply finite_valid_trace_init_to_forget_last in Htr.
      eexists is, tr, _; split; [exact Htr|reflexivity].
    Qed.

    (** Any trace with the 'finite_valid_trace_from' property can be completed
    (to the left) to start in an initial state*)
    Lemma finite_valid_trace_from_complete_left
      (s : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from s tr)
      : exists (is : state) (trs : list transition_item),
        finite_valid_trace is (trs ++ tr) /\
        finite_trace_last is trs = s.
    Proof.
      apply finite_valid_trace_first_pstate in Htr as Hs.
      apply valid_state_has_trace in Hs.
      destruct Hs as [is [trs [Htrs His]]].
      exists is, trs.
      apply finite_valid_trace_from_to_last in Htrs as Hlast.
      rewrite <- Hlast in Htr.
      apply finite_valid_trace_from_to_forget_last in Htrs.
      repeat (split || assumption ||
      apply finite_valid_trace_from_app_iff).
    Qed.

    (** Any trace with the 'finite_valid_trace_from_to' property can be completed
    (to the left) to start in an initial state*)
    Lemma finite_valid_trace_from_to_complete_left
      (s f : state)
      (tr : list transition_item)
      (Htr : finite_valid_trace_from_to s f tr)
      : exists (is : state) (trs : list transition_item),
        finite_valid_trace_init_to is f (trs ++ tr) /\
        finite_trace_last is trs = s.
    Proof.
      assert (valid_state_prop s) as Hs
        by (apply finite_valid_trace_from_to_forget_last,
            finite_valid_trace_first_pstate in Htr; assumption).
      apply valid_state_has_trace in Hs.
      destruct Hs as [is [trs [Htrs His]]].
      exists is, trs.
      split.
      - split;[|assumption].
        apply finite_valid_trace_from_to_app with s;assumption.
      - apply finite_valid_trace_from_to_last in Htrs;assumption.
    Qed.

(** Another benefit of defining traces is that we can succintly
describe indirect transitions between arbitrary pairs of states.

We say that state <<second>> is in state <<first>>'s futures if
there exists a finite (possibly empty) valid trace that begins
with <<first>> and ends in <<second>>.

This relation is often used in stating safety and liveness properties.*)

    Definition in_futures
      (first second : state)
      : Prop :=
      exists (tr : list transition_item),
        finite_valid_trace_from_to first second tr.

    Lemma in_futures_preserving
      (R : state -> state -> Prop)
      (Hpre : PreOrder R)
      (Ht : input_valid_transition_preserving R)
      (s1 s2 : state)
      (Hin : in_futures s1 s2)
      : R s1 s2.
    Proof.
      unfold in_futures in Hin.
      destruct Hin as [tr Htr].
      induction Htr.
      - reflexivity.
      - apply Ht in Ht0.
        transitivity s;assumption.
    Qed.

    Instance eq_equiv : @Equivalence state eq := _.

    Lemma in_futures_strict_preserving
      (R : state -> state -> Prop)
      (Hpre : StrictOrder R)
      (Ht : input_valid_transition_preserving R)
      (s1 s2 : state)
      (Hin : in_futures s1 s2)
      (Hneq : s1 <> s2)
      : R s1 s2.
    Proof.
      apply (StrictOrder_PreOrder eq_equiv) in Hpre.
      - specialize (in_futures_preserving (relation_disjunction R eq) Hpre) as Hpreserve.
        spec Hpreserve.
        + intro; intros. left. apply (Ht s3 s4 l0 om1 om2 Hvalid_transition).
        + spec Hpreserve s1 s2 Hin. destruct Hpreserve; try assumption.
          elim Hneq. assumption.
      - intros x1 x2 Heq. subst. intros y1 y2 Heq. subst.
        split; intro; assumption.
    Qed.

    Lemma in_futures_valid_fst
      (first second : state)
      (Hfuture: in_futures first second)
      : valid_state_prop first.
    Proof.
      destruct Hfuture as [tr Htr].
      apply finite_valid_trace_from_to_forget_last in Htr.
      apply finite_valid_trace_first_pstate in Htr.
      assumption.
    Qed.

    (* begin hide *)

    Lemma in_futures_refl
      (first: state)
      (Hps : valid_state_prop first)
      : in_futures first first.

    Proof.
      exists [].
      constructor.
      assumption.
    Qed.

    Lemma in_futures_trans
      (first second third : state)
      (H12: in_futures first second)
      (H23 : in_futures second third)
      : in_futures first third.
    Proof.
      destruct H12 as [tr12 Htr12].
      destruct H23 as [tr23 Htr23].
      exists (tr12 ++ tr23).
      apply finite_valid_trace_from_to_app with second;assumption.
    Qed.

    Lemma input_valid_transition_in_futures {l s im s' om}
      (Ht : input_valid_transition l (s, im) (s', om))
      : in_futures s s'.
    Proof.
      apply finite_valid_trace_singleton in Ht.
      apply finite_valid_trace_from_add_last with (f := s') in Ht; [|reflexivity].
      eexists. exact Ht.
    Qed.

    Lemma elem_of_trace_in_futures_left is s tr
      (Htr : finite_valid_trace_from_to is s tr)
      : forall item, item ∈ tr -> in_futures (destination item) s.
    Proof.
      intros item Hitem.
      apply elem_of_list_split in Hitem as (pre & suf & Heqtr).
      exists suf.
      replace (destination item)
         with (finite_trace_last is (pre ++ [item]))
           by apply finite_trace_last_is_last.
      eapply finite_valid_trace_from_to_app_split.
      rewrite <- app_assoc. simpl. rewrite <- Heqtr.
      assumption.
    Qed.

    Lemma elem_of_trace_in_futures_right is s tr
      (Htr : finite_valid_trace_from_to is s tr)
      : forall item, item ∈ tr -> in_futures is (destination item).
    Proof.
      intros item Hitem.
      apply elem_of_list_split in Hitem as (pre & suf & Heqtr).
      exists (pre ++ [item]).
      replace (destination item)
         with (finite_trace_last is (pre ++ [item]))
           by apply finite_trace_last_is_last.
      eapply finite_valid_trace_from_to_app_split.
      rewrite <- app_assoc. simpl. rewrite <- Heqtr.
      eassumption.
    Qed.

    Lemma in_futures_witness
      (first second : state)
      (Hfutures : in_futures first second)
      : exists (tr : valid_trace) (n1 n2 : nat),
        n1 <= n2
        /\ trace_nth (proj1_sig tr) n1 = Some first
        /\ trace_nth (proj1_sig tr) n2 = Some second.
    Proof.
      specialize (in_futures_valid_fst first second Hfutures); intro Hps.
      apply valid_state_has_trace in Hps.
      destruct Hps as [prefix_start [prefix_tr [Hprefix_tr Hinit]]].
      destruct Hfutures as [suffix_tr Hsuffix_tr].
      specialize (finite_valid_trace_from_to_app _ _ _ _ _ Hprefix_tr Hsuffix_tr) as Happ.
      apply finite_valid_trace_from_to_forget_last in Happ.
      assert (Htr : valid_trace_prop (Finite prefix_start (prefix_tr ++ suffix_tr)))
        by (split;assumption).
      exists (exist _ _ Htr).
      simpl.
      exists (length prefix_tr), (length prefix_tr + length suffix_tr).
      split;[lia|].
      apply finite_valid_trace_from_to_last in Hprefix_tr.
      apply finite_valid_trace_from_to_last in Hsuffix_tr.
      split.
      - rewrite finite_trace_nth_app1;[|lia].
        rewrite finite_trace_nth_last.
        congruence.
      - rewrite finite_trace_nth_app2;[|lia].
        rewrite Minus.minus_plus.
        rewrite finite_trace_nth_last.
        congruence.
    Qed.

    Definition trace_segment
      (tr : Trace)
      (n1 n2 : nat)
      : list transition_item
      := match tr with
      | Finite s l => list_segment l n1 n2
      | Infinite s l => stream_segment l n1 n2
      end.

    Lemma valid_trace_segment
      (tr : Trace)
      (Htr : valid_trace_prop tr)
      (n1 n2 : nat)
      (Hle : n1 <= n2)
      (first : state)
      (Hfirst : trace_nth tr n1 = Some first)
      : finite_valid_trace_from first (trace_segment tr n1 n2).
    Proof.
      destruct tr as [s tr | s tr]; simpl in *; destruct Htr as [Htr Hinit].
      - apply finite_valid_trace_from_segment with s; try assumption.
      - inversion Hfirst; subst; clear Hfirst.
        apply (infinite_valid_trace_from_segment s tr Htr n1 n2 Hle).
    Qed.

    Inductive Trace_messages : Type :=
    | Finite_messages : list (option message) -> Trace_messages
    | Infinite_messages : Stream (option message) -> Trace_messages.

    Definition protocol_output_messages_trace (tr : valid_trace) : Trace_messages :=
      match proj1_sig tr with
      | Finite _ ls => Finite_messages (List.map output ls)
      | Infinite _ st => Infinite_messages (map output st) end.

    Definition protocol_input_messages_trace (tr : valid_trace) : Trace_messages :=
      match proj1_sig tr with
      | Finite _ ls => Finite_messages (List.map input ls)
      | Infinite _ st => Infinite_messages (map input st) end.

    Definition trace_prefix
               (tr : Trace)
               (last : transition_item)
               (prefix : list transition_item)
      :=
        match tr with
        | Finite s ls => exists suffix, ls = prefix ++ (last :: suffix)
        | Infinite s st => exists suffix, st = stream_app prefix (Cons last suffix)
        end.

    Definition trace_prefix_fn
      (tr : Trace)
      (n : nat)
      : Trace
      :=
      match tr with
      | Finite s ls => Finite s (list_prefix ls n)
      | Infinite s st => Finite s (stream_prefix st n)
      end.

    Lemma trace_prefix_valid
          (tr : valid_trace)
          (last : transition_item)
          (prefix : list transition_item)
          (Hprefix : trace_prefix (proj1_sig tr) last prefix)
      : valid_trace_prop (Finite (trace_first (proj1_sig tr)) (prefix ++ [last])).
    Proof.
      destruct tr as [tr Htr]. simpl in *.
      generalize dependent tr. generalize dependent last.
      apply (rev_ind (fun prefix => forall (last : transition_item) (tr : Trace), valid_trace_prop tr -> trace_prefix tr last prefix -> finite_valid_trace (trace_first tr) (prefix ++ [last]))).
      - intros last tr Htr Hprefix; destruct tr as [ | ]; unfold trace_prefix in Hprefix;   simpl in Hprefix
        ; destruct Hprefix as [suffix Heq]; subst; destruct Htr as [Htr Hinit]
        ; unfold trace_first; simpl; constructor; try assumption
        ; inversion Htr; subst; clear Htr
        ; apply finite_valid_trace_singleton; assumption.
      - intros last_p p Hind last tr Htr Hprefix.
        specialize (Hind last_p tr Htr).
        destruct tr as [ | ]; unfold trace_prefix in Hprefix;   simpl in Hprefix
        ; destruct Hprefix as [suffix Heq]; subst; destruct Htr as [Htr Hinit]; simpl; simpl in Hind
        ; split; try assumption
        .
        + assert
            (Hex : exists suffix0 : list transition_item,
                (p ++ [last_p]) ++ last :: suffix = p ++ last_p :: suffix0
            ) by (exists (last :: suffix); rewrite <- app_assoc; reflexivity)
          ; specialize (Hind Hex); clear Hex
          ; destruct Hind as [Hptr _]
          ; destruct last
          ; apply extend_right_finite_trace_from
          ; try assumption
          .
          rewrite <- (app_cons {| l := l0; input := input0; destination := destination0; output := output0 |} suffix) in Htr.
          rewrite app_assoc in Htr.
          rewrite <- (app_assoc p _ _) in Htr. simpl in Htr.
          rewrite <- app_assoc in Htr.
          specialize
            (finite_valid_trace_consecutive_valid_transition _ _ _ _ _ _ Htr eq_refl).
          simpl.
          rewrite finite_trace_last_is_last. trivial.
        + assert
            (Hex : exists suffix0 : Stream transition_item,
                stream_app (p ++ [last_p])  (Cons last suffix) = stream_app p (Cons last_p suffix0)
            ) by (exists (Cons last suffix); rewrite <- stream_app_assoc; reflexivity)
          ; specialize (Hind Hex); clear Hex
          ; destruct Hind as [Hptr _]
          ; destruct last
          ; apply extend_right_finite_trace_from
          ; try assumption
          .
          rewrite <- stream_app_cons in Htr.
          rewrite stream_app_assoc in Htr.
          rewrite <- (app_assoc p _ _) in Htr. simpl in Htr.
          specialize
            (infinite_valid_trace_consecutive_valid_transition
               s
               (stream_app (p ++ [last_p; {| l := l0; input := input0; destination := destination0; output := output0 |}]) suffix)
               suffix
               p
               last_p
               {| l := l0; input := input0; destination := destination0; output := output0 |}
               Htr
               eq_refl
            ).
          simpl.
          rewrite finite_trace_last_is_last. trivial.
    Qed.


    Definition build_trace_prefix_valid
          {tr : valid_trace}
          {last : transition_item}
          {prefix : list transition_item}
          (Hprefix : trace_prefix (proj1_sig tr) last prefix)
          : valid_trace
      := exist _ (Finite (trace_first (proj1_sig tr)) (prefix ++ [last]))
               (trace_prefix_valid tr last prefix Hprefix).

    Lemma trace_prefix_fn_valid
          (tr : Trace)
          (Htr : valid_trace_prop tr)
          (n : nat)
      : valid_trace_prop (trace_prefix_fn tr n).
    Proof.
      specialize (trace_prefix_valid (exist _ tr Htr)); simpl; intro Hpref.
      remember (trace_prefix_fn tr n) as pref_tr.
      destruct pref_tr as [s l | s l].
      - destruct l as [| item l].
        + destruct tr as [s' l' | s' l']
          ; destruct Htr as [Htr Hinit]
          ; inversion Heqpref_tr; subst
          ; (split;[|assumption])
          ; constructor
          ;  apply initial_state_is_valid;assumption.
        + assert (Hnnil : item ::l <> [])
            by (intro Hnil; inversion Hnil).
          specialize (exists_last Hnnil); intros [prefix [last Heq]].
          rewrite Heq in *; clear Hnnil Heq l item.
          replace s with (trace_first (proj1_sig (exist _ tr Htr)))
          ; try (destruct tr; inversion Heqpref_tr; subst; reflexivity).
          apply trace_prefix_valid.
          remember (prefix ++ [last]) as prefix_last. revert Heqprefix_last.
          destruct tr as [s' l' | s' l']
          ; inversion Heqpref_tr
          ; subst
          ; clear Heqpref_tr
          ; simpl
          ; intro Heqprefix.
          * specialize (list_prefix_suffix l' n); intro Hl'.
            rewrite <- Hl'. rewrite Heqprefix.
            exists (list_suffix l' n).
            rewrite <- app_assoc.
            reflexivity.
          * specialize (stream_prefix_suffix l' n); intro Hl'.
            rewrite <- Hl'. rewrite Heqprefix.
            exists (stream_suffix l' n).
            rewrite <- stream_app_assoc.
            reflexivity.
      - destruct tr as [s' l' | s' l']; inversion Heqpref_tr.
    Qed.

    Lemma valid_trace_nth
      (tr : Trace)
      (Htr : valid_trace_prop tr)
      (n : nat)
      (s : state)
      (Hnth : trace_nth tr n = Some s)
      : valid_state_prop s.
    Proof.
      destruct tr as [s0 l | s0 l]; destruct Htr as [Htr Hinit].
      - specialize (finite_valid_trace_from_suffix s0 l Htr n s Hnth).
        intro Hsuf.
        apply finite_valid_trace_first_pstate in Hsuf.
        assumption.
      - assert (Hle : n <= n) by lia.
        specialize (infinite_valid_trace_from_segment s0 l Htr n n Hle)
        ; simpl; intros Hseg.
        inversion Hnth.
        apply finite_valid_trace_first_pstate in Hseg.
        assumption.
    Qed.

    Lemma in_futures_valid_snd
      (first second : state)
      (Hfutures: in_futures first second)
      : valid_state_prop second.
    Proof.
      specialize (in_futures_witness first second Hfutures)
      ; intros [tr [n1 [n2 [Hle [Hn1 Hn2]]]]].
      destruct tr as [tr Htr]; simpl in Hn2.
      apply valid_trace_nth with tr n2; assumption.
    Qed.

    Lemma in_futures_witness_reverse
      (first second : state)
      (tr : valid_trace)
      (n1 n2 : nat)
      (Hle : n1 <= n2)
      (Hs1 : trace_nth (proj1_sig tr) n1 = Some first)
      (Hs2 : trace_nth (proj1_sig tr) n2 = Some second)
      : in_futures first second.
    Proof.
      destruct tr as [tr Htr].
      simpl in *.
      inversion Hle; subst; clear Hle.
      - rewrite Hs1 in Hs2. inversion Hs2; subst; clear Hs2.
        exists [].
        constructor. apply valid_trace_nth with tr n2; assumption.
      - exists (trace_segment tr n1 (S m)).
        apply finite_valid_trace_from_add_last.
        + apply valid_trace_segment; try assumption. lia.
        + { destruct tr as [s tr | s tr]; simpl.
          - simpl in Hs1, Hs2.
            unfold list_segment.
            rewrite finite_trace_last_suffix.
            apply finite_trace_last_prefix. assumption.
            rewrite list_prefix_length. lia.
            apply finite_trace_nth_length in Hs2. lia.
          - unfold stream_segment.
            rewrite unlock_finite_trace_last.
            rewrite list_suffix_map, stream_prefix_map.
            simpl in Hs2.
            rewrite list_suffix_last.
            + symmetry. rewrite stream_prefix_nth_last.
              unfold Str_nth in Hs2. simpl in Hs2.
              inversion Hs2; subst.
              reflexivity.
            + specialize (stream_prefix_length (Streams.map destination tr) (S m)); intro Hpref_len.
              rewrite Hpref_len.
              lia.
          }
    Qed.
    (* end hide *)

(**
Stating livness properties will require quantifying over complete
executions of the protocol. To make this possible, we will now define
_complete_ [valid_trace]s.

A [valid_trace] is _terminating_ if there's no other [valid_trace]
that contains it as a prefix.
*)

    Definition terminating_trace_prop (tr : Trace) : Prop
       :=
         match tr with
         | Finite s ls =>
             (exists (tr : valid_trace)
             (last : transition_item),
             trace_prefix (proj1_sig tr) last ls) -> False
         | Infinite s ls => False
         end.

(** A [valid_trace] is _complete_, if it is either _terminating_ or infinite.
*)

    Definition complete_trace_prop (tr : Trace) : Prop
       := valid_trace_prop tr
          /\
          match tr with
          | Finite _ _ => terminating_trace_prop tr
          | Infinite _ _ => True
          end.

    (* begin hide *)

    (* Implicitly, the state itself must be in the trace, and minimally the last element of the trace *)
    (* Also implicitly, the trace leading up to the state is finite *)
    (* Defining equivocation on these trace definitions *)

    (* Section 7 :
       A message m received by a valid state s with a transition label l in a
       valid execution trace is called "an equivocation" if it wasn't produced
       in that trace
    *)

    (* 6.2.2 Equivocation-free as a composition constraint *)
    Definition composition_constraint : Type :=
      label -> state * option message -> Prop.

    (* Decidable VLSMs *)

    Class VLSM_vdecidable :=
      { valid_decidable : forall l som, {valid l som} + {~valid l som}
      }.
(* end hide *)
End VLSM.

(** Make all arguments of [valid_state_prop_ind] explicit
    so it will work with the <<induction using>> tactic.
    (closing the section added <<{message}>> as an implicit argument)
 *)
Arguments valid_state_message_prop_ind : clear implicits.
Arguments valid_state_prop_ind : clear implicits.
Arguments finite_valid_trace_from_to_ind : clear implicits.

Arguments finite_valid_trace_rev_ind : clear implicits.
Arguments finite_valid_trace_from_rev_ind : clear implicits.
Arguments finite_valid_trace_from_to_rev_ind : clear implicits.
Arguments finite_valid_trace_init_to_rev_ind : clear implicits.
Arguments finite_valid_trace_init_to_rev_strong_ind : clear implicits.

Arguments extend_right_finite_trace_from [message] (X) [s1] [ts] (Ht12) [l3] [iom3] [s3] [oom3] (Hv23).
Arguments extend_right_finite_trace_from_to [message] (X) [s1] [s2] [ts] (Ht12) [l3] [iom3] [s3] [oom3] (Hv23).

Class TraceWithLast
      (base_prop : forall {message} (X: VLSM message),
      @state _ (@type _ X) -> list transition_item -> Prop)
      (trace_prop : forall {message} (X: VLSM message),
        state -> state -> list transition_item -> Prop) :=
  {valid_trace_add_last: forall [msg] [X: VLSM msg] [s f tr],
     base_prop X s tr -> finite_trace_last s tr = f -> trace_prop X s f tr;
   valid_trace_get_last: forall [msg] [X: VLSM msg] [s f tr],
     trace_prop X s f tr -> finite_trace_last s tr = f;
   valid_trace_last_pstate: forall [msg] [X: VLSM msg] [s f tr],
     trace_prop X s f tr -> valid_state_prop X f;
   valid_trace_forget_last: forall [msg] [X: VLSM msg] [s f tr],
     trace_prop X s f tr -> base_prop X s tr
  }.
Global Hint Mode TraceWithLast - ! : typeclass_instances.
Global Hint Mode TraceWithLast ! - : typeclass_instances.

Definition valid_trace_add_default_last
  `{TraceWithLast base_prop trace_prop}
  [msg] [X:VLSM msg] [s tr] (Htr: base_prop msg X s tr):
    trace_prop msg X s (finite_trace_last s tr) tr.
Proof.
  apply valid_trace_add_last. assumption. reflexivity.
Defined.

Instance trace_with_last_valid_trace_from:
  TraceWithLast (@finite_valid_trace_from) (@finite_valid_trace_from_to)
  := {valid_trace_add_last := @finite_valid_trace_from_add_last;
      valid_trace_get_last := @finite_valid_trace_from_to_last;
      valid_trace_last_pstate := @finite_valid_trace_from_to_last_pstate;
      valid_trace_forget_last := @finite_valid_trace_from_to_forget_last;
     }.

Instance trace_with_last_valid_trace_init:
  TraceWithLast (@finite_valid_trace) (@finite_valid_trace_init_to)
  := {valid_trace_add_last := @finite_valid_trace_init_add_last;
      valid_trace_get_last := @finite_valid_trace_init_to_last;
      valid_trace_last_pstate _ _ _ _ _ H := valid_trace_last_pstate (proj1 H);
      valid_trace_forget_last := @finite_valid_trace_init_to_forget_last;
     }.

Class TraceWithStart
     {message} {X : VLSM message}
     (start : @state message (type X))
     (trace_prop : list (transition_item (type X)) -> Prop) :=
 {valid_trace_first_pstate:
    forall [tr], trace_prop tr -> valid_state_prop X start
 }.
Global Hint Mode TraceWithStart - - - ! : typeclass_instances.

Instance trace_with_start_valid_trace_from message (X: VLSM message) s:
  TraceWithStart s (finite_valid_trace_from X s)
  := {valid_trace_first_pstate := finite_valid_trace_first_pstate X s}.
Instance trace_with_start_valid_trace message (X: VLSM message) s:
  TraceWithStart s (finite_valid_trace X s)
  := {valid_trace_first_pstate tr H := valid_trace_first_pstate (proj1 H)}.
Instance trace_with_start_valid_trace_from_to message (X: VLSM message) s f:
  TraceWithStart s (finite_valid_trace_from_to X s f)
  := {valid_trace_first_pstate tr H := valid_trace_first_pstate (valid_trace_forget_last H)}.
Instance trace_with_start_valid_trace_init_to message (X: VLSM message) s f:
  TraceWithStart s (finite_valid_trace_init_to X s f)
  := {valid_trace_first_pstate tr H := valid_trace_first_pstate (valid_trace_forget_last H)}.

(** *** Pre-loaded VLSMs

Given a VLSM <<X>>, we introduce the _pre-loaded_ version of it,
which is identical to <<X>>, except that it is endowed with the
whole message universe as its initial messages. The high degree
of freedom allowed to the _pre-loaded_ version lets it experience
everything experienced by <<X>> but also other types of behaviour,
including _Byzantine_ behaviour, which makes it a useful concept in
Byzantine fault tolerance analysis.
*)


  Section pre_loaded_with_all_messages_vlsm.
    Context
      {message : Type}
      (X : VLSM message)
      .

  Definition pre_loaded_with_all_messages_vlsm_sig
    : VLSMSign (type X)
    :=
    {| initial_state_prop := vinitial_state_prop X
     ; initial_message_prop := fun message => True
     ; s0 := @s0 _ _ (sign X)
    |}.

  Definition pre_loaded_with_all_messages_vlsm_machine
    : VLSMClass pre_loaded_with_all_messages_vlsm_sig
    :=
    {| transition := vtransition X
     ; valid := vvalid X
    |}.

  Definition pre_loaded_with_all_messages_vlsm
    : VLSM message
    := mk_vlsm pre_loaded_with_all_messages_vlsm_machine.

  (**
    A message which can be emitted during a protocol run of
    the [pre_loaded_with_all_messages_vlsm] is called a [byzantine_message], because
    as shown by Lemmas [byzantine_pre_loaded_with_all_messages] and [pre_loaded_with_all_messages_alt_eq],
    byzantine traces for a [VLSM] are precisely the valid traces
    of the [pre_loaded_with_all_messages_vlsm], hence a byzantine message is any message
    which a byzantine trace [can_emit].
  *)

  Definition byzantine_message_prop
    (m : message)
    : Prop
    := can_emit pre_loaded_with_all_messages_vlsm m.

  Definition byzantine_message : Type
    := sig byzantine_message_prop.

  (* begin hide *)
  Lemma pre_loaded_with_all_messages_message_valid_initial_state_message
    (om : option message)
    : valid_state_message_prop pre_loaded_with_all_messages_vlsm (proj1_sig (vs0 X)) om.
  Proof.
    apply valid_initial_state_message;[apply proj2_sig|].
    destruct om;exact I.
  Qed.

  Lemma pre_loaded_with_all_messages_valid_state_message_preservation
    (s : state)
    (om : option message)
    (Hps : valid_state_message_prop X s om)
    : valid_state_message_prop pre_loaded_with_all_messages_vlsm s om.
  Proof.
    induction Hps.
    - apply (valid_initial_state_message pre_loaded_with_all_messages_vlsm).
      assumption.
      destruct om;exact I.
    - apply (valid_generated_state_message pre_loaded_with_all_messages_vlsm) with s _om _s om l0; assumption.
  Qed.

  Lemma pre_loaded_with_all_messages_valid_state_prop
    (s : state)
    (Hps : valid_state_prop X s)
    : valid_state_prop pre_loaded_with_all_messages_vlsm s.
  Proof.
    unfold valid_state_prop in *.
    destruct Hps as [om Hprs].
    exists om.
    apply pre_loaded_with_all_messages_valid_state_message_preservation.
    intuition.
  Qed.
  (* end hide *)

  Lemma any_message_is_valid_in_preloaded (om: option message):
    option_valid_message_prop pre_loaded_with_all_messages_vlsm om.
  Proof.
    eexists.
    apply pre_loaded_with_all_messages_message_valid_initial_state_message.
  Qed.

  Inductive preloaded_valid_state_prop : state -> Prop :=
  | preloaded_valid_initial_state
      (s:state)
      (Hs: initial_state_prop (VLSMSign:=pre_loaded_with_all_messages_vlsm_sig) s):
         preloaded_valid_state_prop s
  | preloaded_protocol_generated
      (l : label)
      (s : state)
      (Hps : preloaded_valid_state_prop s)
      (om : option message)
      (Hv : valid (VLSMClass:=pre_loaded_with_all_messages_vlsm_machine) l (s, om))
      s' om'
      (Ht : transition (VLSMClass:=pre_loaded_with_all_messages_vlsm_machine) l (s, om) = (s', om'))
    : preloaded_valid_state_prop s'.

  Lemma preloaded_valid_state_prop_iff s:
    valid_state_prop pre_loaded_with_all_messages_vlsm s
    <-> preloaded_valid_state_prop s.
  Proof.
    split.
    - intros [om Hvalid].
      induction Hvalid.
      + apply preloaded_valid_initial_state.
        assumption.
      + apply preloaded_protocol_generated with l0 s om om';assumption.
    - induction 1.
      + exists None.
        apply valid_initial_state_message;[assumption|exact I].
      + exists om'. destruct IHpreloaded_valid_state_prop as [_om Hs].
        specialize (any_message_is_valid_in_preloaded om) as [_s Hom].
        apply (valid_generated_state_message pre_loaded_with_all_messages_vlsm) with s _om _s om l0;assumption.
  Qed.

  Lemma preloaded_weaken_valid_state_message_prop s om:
    valid_state_message_prop X s om ->
    valid_state_message_prop pre_loaded_with_all_messages_vlsm s om.
  Proof.
    induction 1.
    - refine (valid_initial_state_message pre_loaded_with_all_messages_vlsm s Hs om _).
      destruct om;exact I.
    - exact (valid_generated_state_message pre_loaded_with_all_messages_vlsm
                                _ _ IHvalid_state_message_prop1
                                _ _ IHvalid_state_message_prop2 l0 Hv _ _ Ht).
  Qed.

  Lemma preloaded_weaken_input_valid_transition
        l s om s' om':
    input_valid_transition X l (s,om) (s',om') ->
    input_valid_transition pre_loaded_with_all_messages_vlsm l (s,om) (s',om').
  Proof.
    unfold input_valid_transition.
    intros [[[_om valid_s] [_ Hvalid]] Htrans].
    split;[clear Htrans|assumption].
    split.
    - exists _om.
      apply preloaded_weaken_valid_state_message_prop.
      assumption.
    - clear _om valid_s.
      split.
      + apply any_message_is_valid_in_preloaded.
      + assumption.
  Qed.

  Lemma preloaded_weaken_valid_trace_from s tr
    : finite_valid_trace_from X s tr ->
      finite_valid_trace_from pre_loaded_with_all_messages_vlsm s tr.
  Proof.
    intros H. induction H using finite_valid_trace_from_rev_ind.
    - apply (finite_valid_trace_from_empty pre_loaded_with_all_messages_vlsm).
      destruct H as [om H]. exists om.
      revert H. apply preloaded_weaken_valid_state_message_prop.
    - apply (finite_valid_trace_from_app_iff pre_loaded_with_all_messages_vlsm).
      split; [assumption|].
      apply (finite_valid_trace_singleton pre_loaded_with_all_messages_vlsm).
      revert Hx. apply preloaded_weaken_input_valid_transition.
  Qed.

  Lemma pre_traces_with_valid_inputs_are_valid is s tr
    (Htr : finite_valid_trace_init_to pre_loaded_with_all_messages_vlsm is s tr)
    (Hobs : forall m,
      trace_has_message (field_selector input) m tr ->
      valid_message_prop X m
    )
    : finite_valid_trace_init_to X is s tr.
  Proof.
    revert s Htr Hobs.
    induction tr using rev_ind; intros; split
    ; [|apply Htr| | apply Htr]
    ; destruct Htr as [Htr Hinit].
    - inversion Htr. subst.
      apply (finite_valid_trace_from_to_empty X).
      apply initial_state_is_valid. assumption.
    - apply finite_valid_trace_from_to_last in Htr as Hlst.
      apply finite_valid_trace_from_to_app_split in Htr.
      destruct Htr as [Htr Hx].
      specialize (IHtr _ (conj Htr Hinit)).
      spec IHtr.
      { intros. apply Hobs.
        apply trace_has_message_prefix. assumption.
      }
      apply proj1, finite_valid_trace_from_to_forget_last in IHtr.
      apply finite_valid_trace_from_add_last; [|assumption].
      inversion Hx. subst f tl s'.
      apply (extend_right_finite_trace_from X)
      ; [assumption|].
      destruct Ht as [[_ [_ Hv]] Ht].
      apply finite_valid_trace_last_pstate in IHtr as Hplst.
      repeat split; try assumption.
      destruct iom as [m|]; [|apply option_valid_message_None].
      apply option_valid_message_Some.
      apply Hobs.
      apply Exists_app. right.
      apply Exists_cons. left.
      subst. reflexivity.
  Qed.

End pre_loaded_with_all_messages_vlsm.

Lemma non_empty_valid_trace_from_can_produce
  `(X : VLSM message)
  (s : state)
  (m : message)
  : can_produce X s m
  <-> exists (is : state) (tr : list transition_item) (item : transition_item),
    finite_valid_trace X is tr /\
    last_error tr = Some item /\
    destination item = s /\ output item = Some m.
Proof.
  split.
  - intros [(s', om') [l Hsm]].
    destruct (id Hsm) as [[Hp _] _].
    pose proof (finite_valid_trace_singleton _ Hsm) as Htr.
    apply finite_valid_trace_from_complete_left in Htr.
    destruct  Htr as [is [trs [Htrs _]]].
    exists is.
    match type of Htrs with
    | context [_ ++ [?item]] => remember item as lstitem
    end.
    exists (trs ++ [lstitem]). exists lstitem.
    split; [assumption|].
    split; [apply last_error_is_last|].
    subst lstitem.
    split; reflexivity.
  - intros [is [tr [item [Htr [Hitem [Hs Hm]]]]]].
    destruct_list_last tr tr' item' Heq; [inversion Hitem|].
    clear Heq.
    rewrite last_error_is_last in Hitem. inversion Hitem. clear Hitem. subst item'.
    destruct Htr as [Htr _].
    apply finite_valid_trace_from_app_iff in Htr.
    destruct Htr as [_ Htr].
    inversion Htr. clear Htr. subst. simpl in Hm. subst.
    eexists _, l0. apply Ht.
Qed.

(** *** Properties of provably-equal VLSMs

If we know that two VLSMs are provably equal, we could try rewriting by them.
However, that gets usually quite technical. To go around that, we will prove
that there is a [VLSMProjections.VLSM_full_projection] between them which will
allow trace-based results to be easily moved betweent the two VLSMs.

Below are some preliminary results; the actual projection is given in
[VLSMProjections.same_VLSM_full_projection].
*)
Section same_VLSM.

Context
  {message : Type}
  .

Section definitions.

Context
  [X1 X2 : VLSM message]
  (Heq : X1 = X2)
  .

Definition same_VLSM_label_rew (l1 : vlabel X1) : vlabel X2 :=
  eq_rect X1 _ l1 _ Heq.

Definition same_VLSM_state_rew (s1 : vstate X1) : vstate X2 :=
  eq_rect X1 _ s1 _ Heq.

End definitions.

Context
  (X1 X2 : VLSM message)
  (Heq : X1 = X2)
  .

Lemma same_VLSM_valid_preservation l1 s1 om
  : vvalid X1 l1 (s1, om) ->
    vvalid X2 (same_VLSM_label_rew Heq l1) (same_VLSM_state_rew Heq s1, om).
Proof.
  unfold same_VLSM_label_rew, same_VLSM_state_rew.
  revert l1 s1. rewrite Heq.
  intros. assumption.
Qed.

Lemma same_VLSM_transition_preservation l1 s1 om s1' om'
  : vtransition X1 l1 (s1, om) = (s1', om') ->
    vtransition X2 (same_VLSM_label_rew Heq l1) (same_VLSM_state_rew Heq s1, om) =
      (same_VLSM_state_rew Heq s1', om').
Proof.
  unfold same_VLSM_label_rew, same_VLSM_state_rew.
  revert l1 s1 s1'. rewrite Heq.
  intros. assumption.
Qed.

Lemma same_VLSM_initial_state_preservation s1
  : vinitial_state_prop X1 s1 -> vinitial_state_prop X2 (same_VLSM_state_rew Heq s1).
Proof.
  revert s1. unfold same_VLSM_state_rew. rewrite Heq.
  intros. assumption.
Qed.

Lemma same_VLSM_initial_message_preservation m
  : vinitial_message_prop X1 m -> vinitial_message_prop X2 m.
Proof.
  rewrite Heq. exact id.
Qed.

End same_VLSM.
